(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param579 = (-(!((^((8'haa) * (8'hb7))) * ((+(8'hb7)) & (+(8'hb5))))))
, parameter param580 = param579 )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h6ae):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire0;
  input wire signed [(3'h4):(1'h0)] wire1;
  input wire [(3'h6):(1'h0)] wire2;
  input wire signed [(5'h12):(1'h0)] wire3;
  wire signed [(5'h15):(1'h0)] wire532;
  wire [(4'he):(1'h0)] wire531;
  wire signed [(5'h14):(1'h0)] wire530;
  reg [(4'h8):(1'h0)] reg513 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar512 = (1'h0);
  reg [(5'h10):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg528 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar526 = (1'h0);
  reg [(5'h12):(1'h0)] reg525 = (1'h0);
  reg [(4'h9):(1'h0)] reg524 = (1'h0);
  reg [(4'hc):(1'h0)] reg523 = (1'h0);
  reg [(4'hf):(1'h0)] forvar522 = (1'h0);
  reg [(3'h4):(1'h0)] reg521 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg520 = (1'h0);
  reg [(4'hc):(1'h0)] reg519 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar517 = (1'h0);
  reg [(4'hd):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg515 = (1'h0);
  reg [(4'h8):(1'h0)] reg514 = (1'h0);
  reg [(5'h10):(1'h0)] forvar513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg512 = (1'h0);
  reg [(5'h15):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg511 = (1'h0);
  reg [(5'h10):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg507 = (1'h0);
  reg [(4'h8):(1'h0)] reg506 = (1'h0);
  reg signed [(4'he):(1'h0)] reg505 = (1'h0);
  reg [(4'ha):(1'h0)] reg504 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg503 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg502 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar501 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg500 = (1'h0);
  reg [(4'he):(1'h0)] reg499 = (1'h0);
  reg [(4'h8):(1'h0)] reg498 = (1'h0);
  reg [(2'h2):(1'h0)] forvar497 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg496 = (1'h0);
  reg [(3'h6):(1'h0)] forvar490 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg495 = (1'h0);
  reg [(2'h3):(1'h0)] reg494 = (1'h0);
  reg [(5'h12):(1'h0)] reg493 = (1'h0);
  reg [(5'h15):(1'h0)] reg492 = (1'h0);
  reg [(5'h12):(1'h0)] reg491 = (1'h0);
  reg [(4'hf):(1'h0)] reg490 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg489 = (1'h0);
  reg [(4'h8):(1'h0)] reg488 = (1'h0);
  reg [(3'h4):(1'h0)] reg487 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg486 = (1'h0);
  reg [(4'hc):(1'h0)] forvar485 = (1'h0);
  reg [(3'h6):(1'h0)] reg484 = (1'h0);
  reg [(4'hc):(1'h0)] reg483 = (1'h0);
  reg [(4'he):(1'h0)] reg482 = (1'h0);
  reg [(4'hf):(1'h0)] forvar481 = (1'h0);
  reg [(4'hb):(1'h0)] reg480 = (1'h0);
  reg [(5'h10):(1'h0)] reg479 = (1'h0);
  reg [(5'h10):(1'h0)] forvar478 = (1'h0);
  reg [(3'h4):(1'h0)] reg477 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg [(2'h3):(1'h0)] reg474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg473 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar471 = (1'h0);
  reg [(3'h5):(1'h0)] forvar470 = (1'h0);
  wire [(3'h7):(1'h0)] wire469;
  wire signed [(3'h7):(1'h0)] wire468;
  wire [(4'hd):(1'h0)] wire466;
  reg [(4'h9):(1'h0)] forvar4 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5 = (1'h0);
  reg [(4'hd):(1'h0)] reg6 = (1'h0);
  reg [(5'h14):(1'h0)] reg7 = (1'h0);
  reg [(5'h11):(1'h0)] reg8 = (1'h0);
  reg [(5'h11):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg10 = (1'h0);
  reg [(5'h13):(1'h0)] forvar11 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg15 = (1'h0);
  reg [(4'h8):(1'h0)] reg16 = (1'h0);
  reg [(4'hf):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar18 = (1'h0);
  reg [(5'h11):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg20 = (1'h0);
  reg [(4'hc):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar13 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire464;
  wire signed [(4'hd):(1'h0)] wire534;
  wire [(4'hf):(1'h0)] wire535;
  reg signed [(5'h14):(1'h0)] forvar537 = (1'h0);
  reg [(5'h14):(1'h0)] forvar538 = (1'h0);
  reg [(5'h13):(1'h0)] reg539 = (1'h0);
  reg [(5'h11):(1'h0)] reg540 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg541 = (1'h0);
  reg [(3'h4):(1'h0)] reg542 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg543 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg544 = (1'h0);
  reg [(4'hd):(1'h0)] reg545 = (1'h0);
  reg [(4'hc):(1'h0)] forvar546 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg548 = (1'h0);
  reg [(5'h10):(1'h0)] reg549 = (1'h0);
  reg [(5'h14):(1'h0)] forvar550 = (1'h0);
  reg [(5'h12):(1'h0)] reg551 = (1'h0);
  reg signed [(4'he):(1'h0)] reg552 = (1'h0);
  reg [(3'h4):(1'h0)] reg553 = (1'h0);
  reg [(5'h12):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg555 = (1'h0);
  reg [(2'h2):(1'h0)] forvar541 = (1'h0);
  reg signed [(4'he):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar557 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar558 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg559 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg560 = (1'h0);
  reg [(5'h15):(1'h0)] reg561 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg562 = (1'h0);
  reg [(5'h13):(1'h0)] reg563 = (1'h0);
  reg [(4'he):(1'h0)] reg564 = (1'h0);
  reg [(5'h12):(1'h0)] reg565 = (1'h0);
  reg [(3'h6):(1'h0)] reg566 = (1'h0);
  reg [(5'h15):(1'h0)] forvar567 = (1'h0);
  reg [(4'h8):(1'h0)] reg568 = (1'h0);
  reg [(3'h5):(1'h0)] reg569 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg571 = (1'h0);
  reg [(3'h4):(1'h0)] reg572 = (1'h0);
  reg [(4'hd):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg574 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg576 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire577;
  assign y = {wire532,
                 wire531,
                 wire530,
                 reg513,
                 forvar512,
                 reg529,
                 reg528,
                 reg527,
                 forvar526,
                 reg525,
                 reg524,
                 reg523,
                 forvar522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 forvar517,
                 reg516,
                 reg515,
                 reg514,
                 forvar513,
                 reg512,
                 reg501,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 reg498,
                 forvar497,
                 reg496,
                 forvar490,
                 reg485,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 forvar485,
                 reg484,
                 reg483,
                 reg482,
                 forvar481,
                 reg480,
                 reg479,
                 forvar478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 forvar471,
                 forvar470,
                 wire469,
                 wire468,
                 wire466,
                 forvar4,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 forvar11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 forvar18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 forvar13,
                 wire464,
                 wire534,
                 wire535,
                 forvar537,
                 forvar538,
                 reg539,
                 reg540,
                 reg541,
                 reg542,
                 reg543,
                 reg544,
                 reg545,
                 forvar546,
                 reg547,
                 reg548,
                 reg549,
                 forvar550,
                 reg551,
                 reg552,
                 reg553,
                 reg554,
                 reg555,
                 forvar541,
                 reg556,
                 forvar557,
                 forvar558,
                 reg559,
                 reg560,
                 reg561,
                 reg562,
                 reg563,
                 reg564,
                 reg565,
                 reg566,
                 forvar567,
                 reg568,
                 reg569,
                 reg570,
                 reg571,
                 reg572,
                 reg573,
                 reg574,
                 reg575,
                 reg576,
                 wire577,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (1'h0)); forvar4 = (forvar4 + (1'h1)))
        begin
          if ($signed(wire1))
            begin
              reg5 = $signed((wire3[(3'h7):(3'h5)] + wire1));
              reg6 <= {(7'h41)};
              reg7 <= wire1[(3'h4):(1'h1)];
            end
          else
            begin
              reg5 = $unsigned(wire3[(5'h10):(4'hf)]);
              reg6 = $unsigned($signed({{reg7[(1'h0):(1'h0)], $unsigned(reg5)},
                  forvar4}));
              reg7 <= forvar4[(2'h3):(1'h1)];
              reg8 = $unsigned((reg5[(3'h7):(3'h4)] ?
                  (~(8'haa)) : (forvar4[(4'h8):(3'h5)] ?
                      (~^wire1) : ("Q1PudY3tHLghhHTR5Ss" != $unsigned(reg7)))));
            end
        end
      reg9 <= $signed($signed("Dtc"));
      reg10 = wire0[(4'hd):(1'h1)];
      if (($unsigned(reg9[(3'h7):(3'h4)]) ? (8'hbc) : reg8))
        begin
          for (forvar11 = (1'h0); (forvar11 < (1'h0)); forvar11 = (forvar11 + (1'h1)))
            begin
              reg12 <= {$unsigned((~|(wire1[(2'h3):(2'h2)] ?
                      (reg5 ? reg5 : reg6) : {reg6, wire0})))};
              reg13 <= $unsigned("fLCDeIRTRMLRUSu");
              reg14 <= ((^~$unsigned($unsigned($signed(reg7)))) * ((+forvar11) ?
                  $signed((8'haf)) : (($unsigned(reg6) ?
                      (wire3 > forvar11) : (forvar11 ?
                          reg12 : forvar11)) + (^~reg5))));
            end
          if (((^($unsigned((&reg13)) >> $signed(wire0))) ?
              {$unsigned({(~forvar4),
                      (reg7 - (8'ha4))})} : $unsigned($signed(reg10[(3'h6):(2'h3)]))))
            begin
              reg15 <= {({reg10[(3'h4):(2'h3)]} ?
                      (($unsigned(reg7) ^ $signed(wire2)) ?
                          wire1[(2'h3):(1'h1)] : $unsigned((reg9 >> (8'ha6)))) : wire1[(3'h4):(2'h3)]),
                  reg6[(4'h8):(3'h6)]};
              reg16 = (~^((reg12 ~^ ((wire2 ?
                  wire1 : reg13) & wire3)) || ($unsigned((!(7'h41))) ?
                  (+(^wire2)) : wire3)));
            end
          else
            begin
              reg15 = (^~($unsigned(reg15[(1'h0):(1'h0)]) < ($unsigned((reg7 < reg13)) ?
                  $signed(wire2) : (reg13[(4'h8):(3'h7)] ? (+reg9) : wire2))));
              reg16 = $unsigned(reg10[(4'ha):(3'h4)]);
              reg17 <= ($signed((reg7[(3'h4):(2'h2)] <= (^reg6))) >= ($unsigned($signed({(8'hbd)})) ?
                  forvar4 : $unsigned($signed(((8'hb2) != wire3)))));
            end
          for (forvar18 = (1'h0); (forvar18 < (2'h3)); forvar18 = (forvar18 + (1'h1)))
            begin
              reg19 = reg7[(4'h9):(1'h0)];
              reg20 <= ($unsigned($unsigned($signed(reg16))) ?
                  (forvar4 >>> $unsigned((-reg17[(3'h4):(2'h3)]))) : ((~{(~^reg10)}) | $unsigned(reg13[(2'h3):(2'h2)])));
              reg21 <= $signed($unsigned($signed(reg20)));
              reg22 <= wire3;
              reg23 <= $signed(($unsigned($unsigned((forvar11 ?
                  wire0 : (8'hb2)))) << reg14));
            end
        end
      else
        begin
          for (forvar11 = (1'h0); (forvar11 < (2'h3)); forvar11 = (forvar11 + (1'h1)))
            begin
              reg12 = reg21;
            end
          for (forvar13 = (1'h0); (forvar13 < (1'h0)); forvar13 = (forvar13 + (1'h1)))
            begin
              reg14 = $signed(({{"lGdK6TbFrE6Cs", wire2},
                  $unsigned((~(8'had)))} | forvar13));
              reg15 <= ($signed(reg22[(4'he):(1'h0)]) < reg7[(5'h10):(4'hc)]);
              reg16 <= {forvar11[(3'h7):(2'h2)], $signed({$unsigned(reg23)})};
            end
          reg17 <= forvar4[(3'h4):(3'h4)];
        end
    end
  module24 modinst465 (.wire27(reg13), .wire26(forvar11), .wire25(wire0), .clk(clk), .wire29(reg7), .wire28(reg8), .y(wire464));
  module33 modinst467 (wire466, clk, wire464, reg17, reg15, forvar11);
  assign wire468 = reg19[(4'hc):(4'hc)];
  assign wire469 = $unsigned(reg15);
  always
    @(posedge clk) begin
      for (forvar470 = (1'h0); (forvar470 < (2'h2)); forvar470 = (forvar470 + (1'h1)))
        begin
          for (forvar471 = (1'h0); (forvar471 < (2'h3)); forvar471 = (forvar471 + (1'h1)))
            begin
              reg472 = $unsigned(({(8'ha1),
                  (8'ha8)} == $unsigned(wire466[(1'h0):(1'h0)])));
              reg473 <= {wire466[(4'h9):(2'h3)],
                  $unsigned($signed($unsigned((reg6 - reg15))))};
              reg474 = forvar18[(4'h8):(3'h7)];
              reg475 <= reg16;
              reg476 <= $unsigned(((($signed(reg21) & {(8'hb8),
                      reg22}) <<< (~|(wire2 ^~ reg14))) ?
                  ({$unsigned(reg8),
                      {reg20}} && (wire2 - reg473)) : ($signed((reg7 ^ reg17)) ~^ $signed({reg472,
                      forvar13}))));
            end
          reg477 <= ((forvar11 & (reg10 ?
              $unsigned((reg474 - (8'hbf))) : wire0[(4'he):(3'h5)])) + $unsigned({reg20,
              forvar4[(1'h1):(1'h1)]}));
          for (forvar478 = (1'h0); (forvar478 < (1'h1)); forvar478 = (forvar478 + (1'h1)))
            begin
              reg479 <= (-wire2[(2'h2):(1'h1)]);
            end
          reg480 <= wire3[(2'h3):(1'h0)];
          for (forvar481 = (1'h0); (forvar481 < (1'h1)); forvar481 = (forvar481 + (1'h1)))
            begin
              reg482 = $signed(((reg8[(1'h1):(1'h0)] ?
                  wire0 : (+reg16)) ~^ "1B3CLADTXbtMzoFiqte"));
              reg483 <= {(8'hb2), (~$signed(reg5[(2'h3):(1'h0)]))};
            end
        end
      reg484 = {((~{$unsigned(reg13)}) ?
              $signed(reg474[(2'h2):(1'h0)]) : (((reg16 ? (8'hb6) : reg14) ?
                      "MDQ" : (^reg19)) ?
                  (^~reg21) : $signed((forvar470 || reg17)))),
          reg474};
      if (reg479[(4'hb):(3'h6)])
        begin
          for (forvar485 = (1'h0); (forvar485 < (1'h0)); forvar485 = (forvar485 + (1'h1)))
            begin
              reg486 = (+wire469[(3'h5):(2'h2)]);
              reg487 <= $signed($signed($signed({$signed(forvar11)})));
              reg488 = $signed(reg486);
            end
          reg489 <= forvar470;
          reg490 = reg479[(3'h5):(3'h5)];
          if (reg10)
            begin
              reg491 = $unsigned(reg16);
              reg492 = (~{(~(8'hb1))});
              reg493 <= wire468;
            end
          else
            begin
              reg491 = reg16;
              reg492 <= (((8'hba) ? reg482 : reg9) < wire469);
              reg493 <= $signed($signed($unsigned({wire2[(3'h6):(2'h2)]})));
              reg494 = (^reg490[(4'ha):(1'h0)]);
              reg495 <= $unsigned(reg480);
            end
        end
      else
        begin
          if ($signed((reg483 ? wire2 : reg489[(4'h8):(3'h6)])))
            begin
              reg485 = {(!(&(!$unsigned(reg22)))),
                  (reg488 ?
                      forvar481[(4'h8):(3'h5)] : ($signed((forvar11 ?
                          wire3 : reg21)) <<< ((reg472 ?
                          (7'h40) : reg477) * ((8'hae) | reg22))))};
              reg486 <= $unsigned(reg489);
              reg487 <= (reg9 ?
                  ((!reg474[(2'h3):(2'h3)]) - $signed($signed({forvar471,
                      (8'ha0)}))) : ({{{reg20},
                          reg479}} <<< {(reg484 >> reg486[(1'h0):(1'h0)]),
                      $signed(forvar470[(1'h1):(1'h0)])}));
              reg488 = $unsigned({forvar18});
              reg489 <= $signed($unsigned((8'h9e)));
            end
          else
            begin
              reg485 <= wire2[(1'h0):(1'h0)];
            end
          for (forvar490 = (1'h0); (forvar490 < (1'h1)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 <= ((reg475 ?
                  $signed((reg473 ?
                      (reg474 <= (8'h9d)) : (~&reg17))) : $unsigned($signed((!wire468)))) <<< (!(wire464 + $unsigned($signed(reg473)))));
              reg492 <= reg479;
              reg493 = (($signed($signed($unsigned(reg483))) ^~ $unsigned(reg14[(2'h2):(1'h0)])) ^ ($unsigned(($unsigned(wire3) ~^ $unsigned(reg19))) ?
                  (7'h44) : forvar470));
              reg494 = (^(|{(^(reg486 ? reg489 : forvar4)),
                  (((8'ha6) ? (8'hbb) : (7'h42)) ?
                      (^reg486) : wire3[(2'h3):(1'h0)])}));
              reg495 = ((wire2[(3'h5):(3'h4)] < {(reg476[(2'h3):(1'h0)] >> $signed(reg492)),
                  $signed($unsigned(forvar485))}) == (8'h9d));
            end
          reg496 <= reg21;
          for (forvar497 = (1'h0); (forvar497 < (1'h1)); forvar497 = (forvar497 + (1'h1)))
            begin
              reg498 <= reg6[(4'hd):(4'h8)];
              reg499 = $signed(($unsigned($signed({forvar13,
                  wire464})) <<< reg495[(1'h0):(1'h0)]));
            end
          reg500 <= forvar497[(1'h0):(1'h0)];
        end
      if (forvar18)
        begin
          for (forvar501 = (1'h0); (forvar501 < (1'h0)); forvar501 = (forvar501 + (1'h1)))
            begin
              reg502 <= $unsigned((reg495 ? "pkergS9dlwa" : reg474));
              reg503 = {reg484[(3'h5):(3'h5)]};
              reg504 <= $unsigned((8'hb8));
              reg505 = reg476[(1'h1):(1'h0)];
              reg506 <= ($unsigned(forvar13) ?
                  $unsigned(((&forvar490[(2'h3):(2'h3)]) ^ (~forvar490))) : ($unsigned(wire469[(3'h5):(3'h4)]) << reg499[(1'h0):(1'h0)]));
            end
          if (forvar11[(4'hd):(1'h0)])
            begin
              reg507 <= (((reg5[(3'h5):(2'h3)] ^ {(wire464 ? reg474 : reg13),
                  ((8'hbf) ^~ reg503)}) == reg505) <<< ((|((forvar470 ?
                      wire2 : reg498) - (reg506 ? reg489 : reg492))) ?
                  (reg22 >>> $signed(reg498[(3'h5):(3'h5)])) : wire3));
              reg508 <= $unsigned(({((reg14 ?
                          wire0 : reg485) != (reg472 < reg14))} ?
                  forvar470[(1'h1):(1'h0)] : ($signed($signed(wire1)) ?
                      {$signed(reg14)} : reg477[(1'h1):(1'h1)])));
              reg509 = ({reg16[(3'h7):(3'h7)]} ?
                  $signed(reg473) : ((wire3[(5'h10):(4'hf)] ?
                          {reg505} : $unsigned((reg495 + reg494))) ?
                      $unsigned(reg494) : reg482));
              reg510 = $unsigned((reg503[(1'h1):(1'h0)] < (reg476[(3'h4):(3'h4)] * (8'hb1))));
            end
          else
            begin
              reg507 = forvar478;
              reg508 = $signed($unsigned(reg509[(4'hb):(1'h0)]));
              reg509 <= $unsigned(reg482);
              reg510 = ((reg479 ?
                      ((~^(reg475 + reg500)) ?
                          reg474[(1'h1):(1'h1)] : (!$signed(reg486))) : (8'hb9)) ?
                  (^({$signed(reg482)} || ($unsigned(reg491) & $unsigned((8'ha7))))) : reg477);
              reg511 <= (reg494[(1'h1):(1'h0)] & reg16);
            end
        end
      else
        begin
          if (($unsigned((^reg506)) >= (^~($signed((~reg9)) ?
              {reg500} : {(reg506 ~^ reg477), (^~reg505)}))))
            begin
              reg501 <= (~$unsigned($signed(reg21)));
            end
          else
            begin
              reg501 <= $signed(reg17[(1'h1):(1'h1)]);
              reg502 <= "6NRAbWgbGK";
              reg503 <= $signed(($unsigned(reg511) >>> $signed((~$signed(forvar481)))));
              reg504 = ($signed($signed($signed($unsigned(reg483)))) ?
                  $signed(((&{(8'hbc)}) ?
                      (~&$signed((8'hab))) : forvar11[(5'h13):(4'hb)])) : forvar478);
              reg505 = reg480[(4'ha):(2'h2)];
            end
        end
      if (({{$unsigned((^(8'hab)))}, (8'hbe)} >>> (!$signed(reg9))))
        begin
          reg512 <= reg486;
          for (forvar513 = (1'h0); (forvar513 < (1'h1)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 = reg495;
              reg515 = (reg494[(1'h1):(1'h1)] & $signed($signed(reg499[(3'h6):(3'h5)])));
              reg516 <= ((8'hb8) ? reg498[(1'h1):(1'h1)] : reg515);
            end
          for (forvar517 = (1'h0); (forvar517 < (2'h2)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 <= (~&reg5[(4'h8):(2'h3)]);
              reg519 <= $unsigned($signed((^reg502[(2'h2):(1'h1)])));
              reg520 <= (^(-((reg17 ? {(8'h9e), (7'h43)} : $signed(reg482)) ?
                  reg501 : (^~$unsigned(reg5)))));
              reg521 = reg19;
            end
          for (forvar522 = (1'h0); (forvar522 < (1'h1)); forvar522 = (forvar522 + (1'h1)))
            begin
              reg523 <= wire0;
              reg524 = {((|reg10) > "3GECVHds9HbZICAJY4oh")};
              reg525 <= (forvar470 << $unsigned((($unsigned((8'hb8)) >> (wire2 <= (8'ha4))) >> reg23[(2'h2):(1'h0)])));
            end
          for (forvar526 = (1'h0); (forvar526 < (1'h1)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg527 = {(^~{reg15, (+(|reg503))}),
                  ($unsigned((~|forvar18[(4'h9):(1'h1)])) << {(8'hbc),
                      $signed(((8'ha6) ~^ reg511))})};
              reg528 <= reg527;
              reg529 <= reg494;
            end
        end
      else
        begin
          for (forvar512 = (1'h0); (forvar512 < (1'h0)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 <= (forvar501 ?
                  reg480[(3'h6):(1'h1)] : (^$signed($unsigned((8'hb7)))));
              reg514 = {(({(|reg515)} >> (~&(reg502 ? reg515 : reg512))) ?
                      ($unsigned((wire469 != reg490)) & (!reg7)) : reg520[(4'h9):(2'h2)])};
              reg515 = (^~(7'h42));
            end
        end
    end
  assign wire530 = (!$signed((((reg483 ? reg10 : reg491) ?
                       (^forvar501) : $signed(reg513)) & reg503[(1'h0):(1'h0)])));
  assign wire531 = ((({(reg515 & forvar481)} ? $unsigned((~^reg492)) : reg509) ?
                           reg485 : reg503[(2'h3):(1'h0)]) ?
                       (((~&{reg474, forvar478}) ?
                           reg509[(4'ha):(4'h9)] : reg510) >= ((&(^~reg5)) ?
                           (reg507 != $signed(reg485)) : {wire1[(1'h1):(1'h1)],
                               forvar11[(4'ha):(4'h8)]})) : ((forvar485[(3'h4):(1'h0)] ?
                           ((reg474 ^~ reg501) ?
                               (!(8'haa)) : $signed(forvar4)) : {(8'hab),
                               (reg484 == forvar490)}) & (8'ha1)));
  module173 modinst533 (.wire178(reg505), .y(wire532), .wire177(reg23), .wire175(reg521), .wire176(reg9), .clk(clk), .wire174(reg483));
  assign wire534 = forvar526[(5'h12):(1'h1)];
  module373 modinst536 (wire535, clk, reg515, forvar522, wire534, forvar517);
  always
    @(posedge clk) begin
      for (forvar537 = (1'h0); (forvar537 < (2'h3)); forvar537 = (forvar537 + (1'h1)))
        begin
          for (forvar538 = (1'h0); (forvar538 < (1'h1)); forvar538 = (forvar538 + (1'h1)))
            begin
              reg539 <= reg475[(2'h2):(2'h2)];
              reg540 = $unsigned({(~wire468), (8'hba)});
            end
        end
      if (reg514[(2'h2):(1'h1)])
        begin
          if ($signed((~^($unsigned(reg498[(3'h6):(1'h1)]) || $unsigned((&(8'hb4)))))))
            begin
              reg541 <= wire535[(3'h6):(3'h6)];
              reg542 = $signed({(reg21 ? reg5 : {forvar11[(2'h3):(2'h3)]})});
              reg543 = forvar517[(4'hf):(4'hd)];
              reg544 <= {$unsigned(($signed((reg21 >> reg500)) ?
                      $unsigned("MIl1s6Shh0bz") : forvar512[(2'h2):(1'h1)]))};
              reg545 <= {reg525};
            end
          else
            begin
              reg541 <= (reg520[(2'h3):(2'h3)] ?
                  {$unsigned($unsigned((reg509 > reg13))),
                      reg514[(4'h8):(2'h2)]} : ($unsigned((~(reg484 ?
                          reg525 : reg529))) ?
                      (8'hab) : $signed({$signed(forvar513)})));
            end
          for (forvar546 = (1'h0); (forvar546 < (3'h4)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 <= (^~(({(reg9 << wire534)} ?
                      $unsigned((8'hbb)) : {(reg515 ? forvar513 : (8'hbf))}) ?
                  $signed(reg489) : $signed((reg500[(5'h13):(4'ha)] ?
                      (-forvar537) : ((8'ha9) >> forvar471)))));
              reg548 = (^(&($unsigned(reg473[(2'h2):(2'h2)]) ?
                  (~$signed(reg19)) : (+(forvar512 ? reg505 : (8'hae))))));
              reg549 <= "yZFe5leHho";
            end
          for (forvar550 = (1'h0); (forvar550 < (3'h4)); forvar550 = (forvar550 + (1'h1)))
            begin
              reg551 = wire2[(3'h6):(3'h4)];
            end
          if (($signed($unsigned(((-forvar4) & $unsigned(reg499)))) ?
              {(reg480 <<< reg542[(2'h3):(1'h1)]),
                  $signed(reg540[(4'hd):(1'h0)])} : (reg16 ?
                  {((reg473 ? reg491 : (8'hbf)) | "ozh14iTKMr6DRCdoWl"),
                      reg514} : ((^$signed(wire532)) - $signed(wire0)))))
            begin
              reg552 = ($signed((~|forvar538)) ?
                  {reg7[(1'h1):(1'h0)],
                      (|reg513)} : {$signed((forvar11 ~^ $signed(forvar4))),
                      $unsigned("QOD21Ru5QXWa676Ez")});
              reg553 = $signed($signed(({$signed(reg501)} || reg482)));
              reg554 = reg549[(4'ha):(2'h2)];
              reg555 = $unsigned(reg506[(4'h8):(3'h5)]);
            end
          else
            begin
              reg552 = (^(^~(~&{$unsigned(reg491)})));
              reg553 <= {$signed(((+(wire468 ^~ reg516)) ?
                      ((7'h40) || (reg477 >= (8'hb0))) : reg482[(4'hd):(4'ha)]))};
              reg554 = $signed(reg495[(1'h1):(1'h0)]);
              reg555 <= ((~|{(|$unsigned(reg13)),
                  $signed((!(8'hac)))}) < forvar478);
            end
        end
      else
        begin
          for (forvar541 = (1'h0); (forvar541 < (3'h4)); forvar541 = (forvar541 + (1'h1)))
            begin
              reg542 = reg6[(3'h4):(1'h0)];
              reg543 <= {reg504};
              reg544 <= "a9WJpug";
            end
          reg545 <= ($unsigned(reg515[(4'hc):(3'h4)]) && $signed((reg486 ?
              $unsigned(forvar478) : (~|{reg529, (8'hbf)}))));
          for (forvar546 = (1'h0); (forvar546 < (1'h0)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 <= ((+wire535) ? reg502[(1'h0):(1'h0)] : "BKQX");
            end
          reg548 = "6ap68qRwNkaZnKmTMwP";
        end
      reg556 = forvar517;
      for (forvar557 = (1'h0); (forvar557 < (2'h2)); forvar557 = (forvar557 + (1'h1)))
        begin
          for (forvar558 = (1'h0); (forvar558 < (2'h3)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 = ($unsigned("") ~^ ((({wire530} ?
                          $signed((8'hb7)) : (reg10 ? wire535 : wire530)) ?
                      {reg529} : forvar550[(3'h5):(1'h1)]) ?
                  (($signed(reg473) ^~ $signed(forvar497)) || ((reg547 ?
                      reg472 : reg23) || reg511)) : (reg513[(2'h3):(2'h2)] ?
                      reg500[(2'h3):(2'h2)] : ($unsigned(forvar485) >>> $unsigned((8'hb5))))));
              reg560 <= $unsigned((!$signed($signed((reg553 - reg8)))));
              reg561 <= (|($signed(($signed(wire535) >> (-forvar497))) ?
                  $signed(reg519) : (-$signed((reg486 > wire464)))));
            end
          if ((^~((reg547 ?
                  ($unsigned(forvar546) <= "4zSWcLt1z34tQS") : $signed($unsigned(reg516))) ?
              (~&($signed(forvar4) ?
                  (|reg494) : reg16)) : (({(8'hb7)} >= (~|reg485)) ?
                  {reg486, reg488} : ($unsigned(forvar471) < (reg472 ?
                      forvar485 : reg504))))))
            begin
              reg562 <= (reg559 ?
                  ($signed($unsigned($signed((8'hbb)))) ~^ $signed($unsigned(reg475))) : ((reg545[(2'h3):(1'h1)] ^~ reg9) == ({(reg22 & reg507)} ?
                      $unsigned(((8'hbe) ? forvar4 : (8'ha9))) : ((forvar18 ?
                              reg529 : wire535) ?
                          reg520[(1'h1):(1'h1)] : $unsigned(reg10)))));
              reg563 <= forvar526;
              reg564 <= (($signed("lqgJ8kUKWpCpiwBhn5ep") ~^ ($unsigned((reg552 ?
                          reg549 : reg540)) ?
                      (forvar538 && $signed(reg514)) : (reg503 ?
                          ((8'ha9) || reg14) : {reg479, forvar546}))) ?
                  reg503 : $unsigned(reg514[(3'h6):(2'h2)]));
              reg565 = $unsigned((reg518 ?
                  reg5[(2'h3):(1'h1)] : wire534[(3'h4):(1'h1)]));
              reg566 = $unsigned($unsigned({(~reg488),
                  forvar557[(3'h6):(2'h2)]}));
            end
          else
            begin
              reg562 = $signed((reg8 >> ($signed(reg16) ^ reg496)));
              reg563 <= (forvar550 < forvar478[(4'hb):(3'h4)]);
            end
          for (forvar567 = (1'h0); (forvar567 < (2'h3)); forvar567 = (forvar567 + (1'h1)))
            begin
              reg568 = $signed((8'hac));
              reg569 = (8'hb5);
              reg570 <= $signed((8'ha4));
              reg571 = (~^((((reg528 ? reg482 : reg496) ?
                      (forvar490 ?
                          wire469 : forvar537) : (forvar512 + reg492)) & (+wire2[(1'h1):(1'h1)])) ?
                  reg515[(3'h4):(1'h1)] : wire532));
            end
          if (forvar490[(3'h5):(3'h5)])
            begin
              reg572 <= forvar541[(1'h0):(1'h0)];
              reg573 = forvar485[(2'h2):(1'h0)];
              reg574 = reg506[(1'h1):(1'h1)];
              reg575 <= (|$unsigned(({reg13, (reg19 >= reg559)} ?
                  $signed({reg505}) : reg524)));
              reg576 <= $unsigned(reg519[(4'ha):(1'h1)]);
            end
          else
            begin
              reg572 = (8'hbf);
              reg573 <= (((reg512 ?
                      forvar558 : ($unsigned(reg560) ^~ (reg562 * reg554))) ?
                  reg552[(3'h4):(2'h2)] : $unsigned(((reg539 ?
                      forvar11 : reg473) | {forvar501,
                      reg479}))) > (&(reg21[(3'h5):(2'h2)] ?
                  {(|(8'hbf))} : reg564)));
              reg574 = ($signed($signed((!reg7[(3'h7):(3'h4)]))) && {forvar470[(1'h1):(1'h1)],
                  forvar471[(3'h5):(3'h4)]});
            end
        end
    end
  module173 modinst578 (wire577, clk, reg495, forvar537, reg8, reg484, reg573);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module24
#( parameter param463 = (((~(-((8'hbf) ? (8'had) : (8'hb6)))) ? {(~|(7'h43))} : ({(~(8'hb1)), ((8'hae) ? (8'hab) : (8'hb1))} ? ((~&(8'hb1)) ? {(8'hb2)} : (8'hae)) : ((&(8'hbc)) ? ((7'h40) ? (8'ha8) : (8'hb3)) : (7'h44)))) >>> ((~^(((7'h42) ? (8'hb0) : (8'hb1)) ? ((8'haa) <<< (7'h42)) : {(8'hba), (8'hac)})) & ((8'hab) ? ((|(8'hb4)) ? ((8'hae) || (8'h9c)) : ((8'ha9) ^ (8'ha0))) : {((7'h44) ? (8'h9d) : (8'hb2))}))) )
(y, clk, wire25, wire26, wire27, wire28, wire29);
  output wire [(32'h364):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire25;
  input wire signed [(5'h13):(1'h0)] wire26;
  input wire [(4'hf):(1'h0)] wire27;
  input wire [(4'hd):(1'h0)] wire28;
  input wire signed [(5'h14):(1'h0)] wire29;
  wire signed [(3'h6):(1'h0)] wire462;
  wire signed [(3'h7):(1'h0)] wire460;
  wire [(4'hf):(1'h0)] wire30;
  wire signed [(3'h7):(1'h0)] wire31;
  wire [(5'h11):(1'h0)] wire32;
  wire signed [(4'h8):(1'h0)] wire99;
  reg [(4'h8):(1'h0)] forvar101 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar102 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg104 = (1'h0);
  reg [(4'hd):(1'h0)] reg105 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg106 = (1'h0);
  reg [(5'h14):(1'h0)] forvar107 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg108 = (1'h0);
  reg [(4'hd):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg110 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg111 = (1'h0);
  reg [(4'h8):(1'h0)] reg112 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar113 = (1'h0);
  reg [(3'h5):(1'h0)] reg114 = (1'h0);
  reg [(5'h11):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg [(5'h11):(1'h0)] forvar118 = (1'h0);
  reg [(2'h3):(1'h0)] forvar119 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg122 = (1'h0);
  reg [(4'hf):(1'h0)] reg123 = (1'h0);
  reg [(4'h8):(1'h0)] forvar124 = (1'h0);
  reg [(4'hb):(1'h0)] reg125 = (1'h0);
  reg [(3'h7):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg127 = (1'h0);
  reg [(5'h14):(1'h0)] reg128 = (1'h0);
  reg [(2'h3):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar130 = (1'h0);
  reg [(4'h9):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg132 = (1'h0);
  reg [(5'h13):(1'h0)] reg133 = (1'h0);
  reg [(3'h6):(1'h0)] reg134 = (1'h0);
  reg [(3'h4):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar136 = (1'h0);
  reg [(4'h8):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg138 = (1'h0);
  reg [(3'h4):(1'h0)] reg139 = (1'h0);
  reg [(4'ha):(1'h0)] reg140 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar141 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(4'he):(1'h0)] reg141 = (1'h0);
  reg [(4'ha):(1'h0)] reg143 = (1'h0);
  reg [(4'hf):(1'h0)] reg144 = (1'h0);
  reg [(5'h15):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar146 = (1'h0);
  reg [(3'h5):(1'h0)] forvar147 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg148 = (1'h0);
  reg [(4'hf):(1'h0)] reg149 = (1'h0);
  reg [(3'h5):(1'h0)] reg150 = (1'h0);
  reg [(2'h2):(1'h0)] reg151 = (1'h0);
  reg [(4'ha):(1'h0)] reg152 = (1'h0);
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  reg [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar156 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg157 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg158 = (1'h0);
  reg [(4'hd):(1'h0)] forvar159 = (1'h0);
  reg [(5'h14):(1'h0)] forvar160 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg161 = (1'h0);
  reg [(4'he):(1'h0)] reg162 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg163 = (1'h0);
  reg [(4'h8):(1'h0)] forvar164 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar165 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg167 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg168 = (1'h0);
  reg [(4'h8):(1'h0)] forvar169 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg170 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire171;
  wire [(5'h14):(1'h0)] wire172;
  wire signed [(3'h5):(1'h0)] wire371;
  assign y = {wire462,
                 wire460,
                 wire30,
                 wire31,
                 wire32,
                 wire99,
                 forvar101,
                 forvar102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 forvar107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 forvar113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 forvar118,
                 forvar119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 forvar124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 reg129,
                 forvar130,
                 reg131,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 forvar136,
                 reg137,
                 reg138,
                 reg139,
                 reg140,
                 forvar141,
                 reg142,
                 reg136,
                 reg141,
                 reg143,
                 reg144,
                 reg145,
                 forvar146,
                 forvar147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 reg152,
                 reg153,
                 reg154,
                 reg155,
                 forvar156,
                 reg157,
                 reg158,
                 forvar159,
                 forvar160,
                 reg161,
                 reg162,
                 reg163,
                 forvar164,
                 forvar165,
                 reg166,
                 reg167,
                 reg168,
                 forvar169,
                 reg170,
                 wire171,
                 wire172,
                 wire371,
                 (1'h0)};
  assign wire30 = $unsigned(($signed($unsigned({wire27})) != ($signed((-wire26)) ?
                      ($signed(wire29) ?
                          wire25[(3'h6):(3'h4)] : ((8'h9e) ?
                              wire29 : wire27)) : wire25[(1'h0):(1'h0)])));
  assign wire31 = $unsigned({$signed(((8'h9e) | wire30))});
  assign wire32 = ((~"7") ? (8'haf) : {wire30, (8'hbd)});
  module33 modinst100 (wire99, clk, wire26, wire30, wire32, wire29);
  always
    @(posedge clk) begin
      for (forvar101 = (1'h0); (forvar101 < (2'h3)); forvar101 = (forvar101 + (1'h1)))
        begin
          for (forvar102 = (1'h0); (forvar102 < (1'h1)); forvar102 = (forvar102 + (1'h1)))
            begin
              reg103 = ((&wire29) ? $signed({wire27}) : $unsigned(wire27));
              reg104 = $signed({wire28, (!{(+wire30), (~reg103)})});
              reg105 <= wire32;
              reg106 <= wire27;
            end
          for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
            begin
              reg108 = {$unsigned(reg104[(3'h5):(1'h0)])};
              reg109 = ($signed((~^((reg108 <<< wire30) ?
                      $unsigned(wire28) : $unsigned((8'had))))) ?
                  reg105 : reg108);
              reg110 <= (!((^~wire28[(4'hd):(2'h3)]) ?
                  ($unsigned($signed(reg103)) != $unsigned((~^reg106))) : $unsigned($unsigned(reg105))));
              reg111 = $unsigned(forvar107);
              reg112 <= $signed("PHbWMl545Sk20xvGC");
            end
          for (forvar113 = (1'h0); (forvar113 < (3'h4)); forvar113 = (forvar113 + (1'h1)))
            begin
              reg114 <= reg104[(3'h6):(1'h0)];
              reg115 = wire32;
              reg116 <= (wire28[(2'h2):(1'h1)] >= $signed(($signed(forvar101) ?
                  (forvar102[(1'h1):(1'h0)] ?
                      $unsigned(wire32) : wire26[(3'h6):(3'h6)]) : (+{forvar107}))));
              reg117 = {$signed($unsigned($signed((wire30 >>> wire32)))),
                  reg112[(1'h1):(1'h0)]};
            end
        end
      for (forvar118 = (1'h0); (forvar118 < (2'h3)); forvar118 = (forvar118 + (1'h1)))
        begin
          for (forvar119 = (1'h0); (forvar119 < (3'h4)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 = reg115;
              reg121 <= ((^(~^(~&(reg108 ?
                  wire31 : wire30)))) ^~ (($unsigned($signed((8'ha2))) << $signed($unsigned(reg116))) + "ZLiLAa1YEyn84anQRg"));
              reg122 = reg121;
              reg123 <= wire26[(4'hd):(4'hc)];
            end
          for (forvar124 = (1'h0); (forvar124 < (3'h4)); forvar124 = (forvar124 + (1'h1)))
            begin
              reg125 <= (-$signed(forvar101[(2'h2):(2'h2)]));
              reg126 <= {$signed(wire29[(2'h2):(2'h2)])};
              reg127 = wire30;
              reg128 <= (($unsigned($unsigned($signed(wire27))) + $signed(($signed(forvar124) ?
                  $signed(reg109) : reg116[(2'h2):(1'h0)]))) & (~&(8'ha2)));
            end
          reg129 <= {wire32[(3'h4):(2'h2)], reg110};
          for (forvar130 = (1'h0); (forvar130 < (3'h4)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= $signed(reg125[(3'h7):(1'h1)]);
              reg132 = $unsigned($signed({reg111[(2'h2):(1'h1)],
                  $signed((8'ha3))}));
              reg133 = wire26;
              reg134 <= $signed(wire29[(5'h10):(3'h7)]);
              reg135 <= (&((forvar101[(2'h2):(1'h1)] * {$unsigned(reg115)}) && {(forvar124 & $signed(reg129)),
                  {$unsigned(wire31), $unsigned(reg111)}}));
            end
        end
      if (reg114[(2'h2):(1'h1)])
        begin
          for (forvar136 = (1'h0); (forvar136 < (2'h2)); forvar136 = (forvar136 + (1'h1)))
            begin
              reg137 = (+$unsigned((^~reg116[(2'h3):(2'h2)])));
              reg138 <= ($unsigned($unsigned($signed(((8'ha6) + reg114)))) <= $unsigned($signed((reg111[(2'h2):(1'h0)] <= (wire31 <= reg127)))));
              reg139 <= (((-(reg103 ?
                      $unsigned(reg120) : (wire32 ? forvar107 : (7'h42)))) ?
                  ($signed((!forvar118)) ?
                      {(^~reg138)} : $signed({reg114,
                          reg109})) : (8'hb9)) >>> reg112);
              reg140 = (8'hb9);
            end
          for (forvar141 = (1'h0); (forvar141 < (3'h4)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg142 <= $signed(reg128);
            end
        end
      else
        begin
          reg136 = $unsigned(forvar113[(4'ha):(2'h2)]);
          reg137 = forvar107[(5'h14):(4'hb)];
          if (wire30[(4'hb):(3'h4)])
            begin
              reg138 <= reg131[(1'h1):(1'h1)];
              reg139 <= $signed(wire30);
            end
          else
            begin
              reg138 <= ({(-reg135[(3'h4):(2'h2)])} < (~|({{reg142},
                  $unsigned(reg133)} >>> ((reg138 ? reg108 : reg127) ?
                  (reg131 ? wire32 : forvar130) : $unsigned(reg110)))));
              reg139 <= $signed({(&reg117[(2'h3):(2'h2)]),
                  $signed(({wire31} >>> reg114))});
              reg140 = ($unsigned(({forvar102[(1'h1):(1'h1)]} ?
                  wire25[(4'ha):(1'h0)] : (^~(reg108 ?
                      wire31 : forvar102)))) && (&(^((reg131 ?
                      wire99 : reg125) ?
                  ((8'hb5) ? wire25 : reg120) : reg126[(1'h0):(1'h0)]))));
              reg141 = (&reg116[(3'h4):(1'h1)]);
            end
        end
      reg143 = $unsigned(reg121[(3'h5):(2'h3)]);
      reg144 <= (reg122 ?
          (!(({wire30, (8'had)} ?
                  $signed((8'h9f)) : ((8'ha9) ? forvar118 : reg121)) ?
              ((7'h44) & (reg111 ?
                  reg137 : forvar102)) : forvar101[(1'h1):(1'h1)])) : $signed((~^((reg121 ?
              wire30 : wire28) - ((8'haf) ^ reg111)))));
    end
  always
    @(posedge clk) begin
      reg145 <= reg141[(4'h9):(4'h9)];
      for (forvar146 = (1'h0); (forvar146 < (2'h2)); forvar146 = (forvar146 + (1'h1)))
        begin
          for (forvar147 = (1'h0); (forvar147 < (1'h1)); forvar147 = (forvar147 + (1'h1)))
            begin
              reg148 <= (7'h42);
              reg149 <= ((("Anhg" ~^ (^~wire32[(4'hf):(1'h0)])) & (-"XgcVPF1YJ3qA0yo8")) ?
                  reg112 : {reg136[(2'h3):(1'h0)]});
            end
          if ((8'hb2))
            begin
              reg150 = (^$unsigned({((~&reg145) ?
                      reg117[(4'ha):(3'h4)] : (forvar146 ? reg112 : (8'ha7))),
                  forvar119[(2'h3):(1'h0)]}));
              reg151 <= ((^~($unsigned($unsigned(forvar130)) >> wire27[(1'h0):(1'h0)])) != $unsigned(reg139[(1'h0):(1'h0)]));
              reg152 = $signed((8'h9f));
            end
          else
            begin
              reg150 <= wire31[(1'h1):(1'h1)];
            end
          if ({$unsigned(($signed($signed((8'hbf))) & $signed($signed(reg104))))})
            begin
              reg153 = $signed(reg125);
            end
          else
            begin
              reg153 = $signed((+($signed($unsigned(wire99)) >> ({reg110} ?
                  (8'h9c) : {forvar147}))));
              reg154 <= reg109[(3'h4):(1'h1)];
              reg155 <= reg145[(4'hb):(2'h3)];
            end
          for (forvar156 = (1'h0); (forvar156 < (3'h4)); forvar156 = (forvar156 + (1'h1)))
            begin
              reg157 <= forvar101[(3'h6):(2'h2)];
            end
          reg158 <= "1iAN2bus6DDExfv7QI0";
        end
      for (forvar159 = (1'h0); (forvar159 < (3'h4)); forvar159 = (forvar159 + (1'h1)))
        begin
          for (forvar160 = (1'h0); (forvar160 < (1'h0)); forvar160 = (forvar160 + (1'h1)))
            begin
              reg161 = wire30[(4'hf):(4'hb)];
              reg162 <= ($unsigned(((reg110[(3'h4):(3'h4)] <<< (reg150 || wire28)) & wire27[(4'ha):(2'h3)])) ?
                  ((^reg106) || wire26[(4'h8):(1'h1)]) : (~&$signed($signed((reg154 ~^ forvar146)))));
              reg163 <= $unsigned(reg151[(1'h0):(1'h0)]);
            end
        end
      for (forvar164 = (1'h0); (forvar164 < (1'h0)); forvar164 = (forvar164 + (1'h1)))
        begin
          for (forvar165 = (1'h0); (forvar165 < (1'h1)); forvar165 = (forvar165 + (1'h1)))
            begin
              reg166 <= ((((^~reg141[(1'h1):(1'h1)]) ?
                  ($unsigned(forvar102) ?
                      reg158[(2'h3):(1'h1)] : wire31) : (|$unsigned((7'h42)))) + $signed($signed(forvar159[(4'h9):(1'h0)]))) ^~ reg142[(3'h5):(1'h1)]);
              reg167 <= wire30;
            end
          reg168 <= ($unsigned(forvar101) ?
              (~&$signed({$unsigned((8'ha0)),
                  reg111[(3'h5):(3'h5)]})) : (~{"NzYqbA", (8'hbb)}));
          for (forvar169 = (1'h0); (forvar169 < (3'h4)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg170 = forvar147;
            end
        end
    end
  assign wire171 = (((~((reg116 ? (8'hbc) : reg104) ^~ $signed(reg161))) ?
                       "" : $unsigned((^~{forvar141,
                           wire30}))) ^~ $signed(((reg136[(2'h3):(1'h1)] != $unsigned(reg158)) ?
                       $unsigned($unsigned(wire25)) : ((reg103 ?
                               reg103 : reg136) ?
                           ((8'hbe) < reg109) : (reg122 ?
                               wire27 : forvar124)))));
  assign wire172 = ((($signed((reg135 ? reg161 : reg123)) ?
                       ({reg145} ? wire171 : forvar124) : $unsigned((reg104 ?
                           reg125 : forvar113))) == (reg167 ~^ wire29)) ^ reg105[(4'hc):(4'h8)]);
  module173 modinst372 (wire371, clk, reg140, reg157, wire172, reg127, forvar136);
  module373 modinst461 (wire460, clk, reg144, reg115, wire25, reg145);
  assign wire462 = (^~($unsigned($signed(reg133[(3'h5):(2'h2)])) ?
                       $signed($unsigned((~&reg155))) : $unsigned((reg139 <<< (reg109 <= forvar146)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module373
#(parameter param459 = (+((!{(~|(8'hbe))}) + (8'hb9))))
(y, clk, wire377, wire376, wire375, wire374);
  output wire [(32'h3ee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire377;
  input wire [(4'hf):(1'h0)] wire376;
  input wire signed [(4'hd):(1'h0)] wire375;
  input wire signed [(5'h15):(1'h0)] wire374;
  reg [(5'h12):(1'h0)] reg458 = (1'h0);
  reg [(5'h14):(1'h0)] reg457 = (1'h0);
  reg [(3'h5):(1'h0)] reg456 = (1'h0);
  reg [(5'h14):(1'h0)] reg455 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg454 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg452 = (1'h0);
  reg [(2'h3):(1'h0)] reg451 = (1'h0);
  reg [(4'he):(1'h0)] reg450 = (1'h0);
  reg [(4'hd):(1'h0)] reg449 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar448 = (1'h0);
  reg [(5'h10):(1'h0)] reg447 = (1'h0);
  reg [(5'h14):(1'h0)] reg446 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar445 = (1'h0);
  reg [(5'h15):(1'h0)] forvar444 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire443;
  reg [(5'h11):(1'h0)] reg442 = (1'h0);
  reg [(4'ha):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg440 = (1'h0);
  reg [(3'h7):(1'h0)] forvar439 = (1'h0);
  reg [(4'hf):(1'h0)] reg438 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar436 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar433 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg435 = (1'h0);
  reg [(4'ha):(1'h0)] reg434 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg431 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg430 = (1'h0);
  reg [(5'h11):(1'h0)] reg429 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg428 = (1'h0);
  reg [(4'he):(1'h0)] forvar427 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar426 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg424 = (1'h0);
  reg [(4'hf):(1'h0)] reg423 = (1'h0);
  reg [(3'h4):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg421 = (1'h0);
  reg [(5'h13):(1'h0)] reg420 = (1'h0);
  reg [(5'h10):(1'h0)] reg419 = (1'h0);
  reg [(3'h7):(1'h0)] forvar418 = (1'h0);
  reg [(5'h15):(1'h0)] reg417 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg416 = (1'h0);
  reg [(4'h9):(1'h0)] forvar415 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg413 = (1'h0);
  reg [(2'h2):(1'h0)] forvar412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg411 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg410 = (1'h0);
  reg [(5'h14):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar408 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg407 = (1'h0);
  reg [(5'h13):(1'h0)] reg406 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg405 = (1'h0);
  reg [(4'hb):(1'h0)] forvar404 = (1'h0);
  reg [(2'h2):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg402 = (1'h0);
  reg [(4'ha):(1'h0)] reg401 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg399 = (1'h0);
  reg [(5'h15):(1'h0)] forvar398 = (1'h0);
  reg [(2'h3):(1'h0)] forvar397 = (1'h0);
  reg [(5'h14):(1'h0)] reg396 = (1'h0);
  reg [(4'ha):(1'h0)] reg395 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg394 = (1'h0);
  reg [(5'h11):(1'h0)] reg393 = (1'h0);
  reg [(5'h15):(1'h0)] reg392 = (1'h0);
  reg [(3'h7):(1'h0)] reg391 = (1'h0);
  reg [(4'h8):(1'h0)] reg390 = (1'h0);
  reg [(2'h2):(1'h0)] reg389 = (1'h0);
  reg [(4'hb):(1'h0)] reg388 = (1'h0);
  reg [(4'he):(1'h0)] reg387 = (1'h0);
  reg [(4'hb):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar384 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg382 = (1'h0);
  reg [(4'hc):(1'h0)] forvar381 = (1'h0);
  reg [(4'hb):(1'h0)] reg380 = (1'h0);
  wire [(5'h11):(1'h0)] wire379;
  wire signed [(4'ha):(1'h0)] wire378;
  assign y = {reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 forvar448,
                 reg447,
                 reg446,
                 forvar445,
                 forvar444,
                 wire443,
                 reg442,
                 reg441,
                 reg440,
                 forvar439,
                 reg438,
                 reg437,
                 forvar436,
                 forvar433,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 forvar418,
                 reg417,
                 reg416,
                 forvar415,
                 reg414,
                 reg413,
                 forvar412,
                 reg411,
                 reg410,
                 reg409,
                 forvar408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 forvar398,
                 forvar397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 forvar384,
                 reg383,
                 reg382,
                 forvar381,
                 reg380,
                 wire379,
                 wire378,
                 (1'h0)};
  assign wire378 = {wire374,
                       ((wire374[(4'hd):(4'h8)] ?
                           {(wire376 & wire375)} : $signed(((7'h44) ?
                               wire375 : (8'ha0)))) << {$unsigned("yIZqTJho7DII"),
                           (7'h43)})};
  assign wire379 = (wire378[(3'h7):(2'h3)] ?
                       "E9XY8GbPS" : (+$signed(wire375[(3'h7):(1'h1)])));
  always
    @(posedge clk) begin
      reg380 = $unsigned(((~wire374) && wire378[(2'h2):(2'h2)]));
      for (forvar381 = (1'h0); (forvar381 < (3'h4)); forvar381 = (forvar381 + (1'h1)))
        begin
          reg382 <= $unsigned({$signed(wire376[(4'he):(4'hd)]),
              {wire375[(3'h7):(3'h5)],
                  $signed((wire375 ? wire379 : wire379))}});
          reg383 = (^reg382);
        end
      for (forvar384 = (1'h0); (forvar384 < (3'h4)); forvar384 = (forvar384 + (1'h1)))
        begin
          reg385 = ($signed((^~wire377[(2'h2):(1'h0)])) <<< (~|(^~$unsigned({wire374,
              forvar381}))));
          if ($unsigned($signed({$unsigned(wire374[(4'hc):(2'h3)]),
              $unsigned((-(7'h42)))})))
            begin
              reg386 = $unsigned($unsigned(wire374));
              reg387 = (wire374 << ({wire379[(4'h9):(3'h4)]} - $signed($signed({(8'ha5)}))));
              reg388 = reg380;
              reg389 <= wire376[(2'h2):(2'h2)];
              reg390 <= $signed(($unsigned($unsigned($unsigned((8'hb8)))) & ((reg383[(1'h1):(1'h1)] ?
                  $signed((8'haf)) : (|forvar381)) << (reg385[(1'h1):(1'h1)] ?
                  (8'ha1) : $signed(reg386)))));
            end
          else
            begin
              reg386 = $signed(($signed((8'hb3)) * (($unsigned(wire376) > $signed((8'ha7))) <<< $unsigned((wire377 ?
                  (8'hb4) : reg386)))));
              reg387 = {($signed((~|$signed(reg380))) ?
                      $signed((~&$unsigned(reg389))) : {$unsigned(wire379)})};
            end
          reg391 = $signed((&wire379));
          if ((((^(8'h9c)) != $unsigned(({wire374, (8'h9e)} ?
                  $signed((8'hb1)) : $signed(wire379)))) ?
              ((|$signed((reg383 ?
                  wire376 : (8'hbf)))) >>> $signed({reg390[(1'h1):(1'h1)]})) : reg380[(4'h8):(2'h2)]))
            begin
              reg392 <= (8'hb5);
            end
          else
            begin
              reg392 <= (+reg389[(1'h1):(1'h1)]);
              reg393 = ($signed((forvar384[(3'h5):(1'h1)] ?
                      "n3Pao2bzppV1KuWKWpE" : $signed($signed(forvar384)))) ?
                  (&({$signed(wire375),
                      wire377[(4'hd):(4'hb)]} << $unsigned($unsigned((8'ha3))))) : (|$unsigned((reg387[(3'h4):(3'h4)] ?
                      ((8'hba) || reg392) : $unsigned(reg387)))));
              reg394 <= ({(~$signed((reg382 & reg382)))} + ((&$signed(wire375)) ?
                  ((!forvar381) ~^ ($unsigned(wire375) ^~ wire378[(3'h6):(1'h0)])) : (~$unsigned((reg387 != reg380)))));
              reg395 <= ((((reg387 ?
                  (wire375 ?
                      reg383 : (8'hb1)) : reg394[(4'ha):(1'h0)]) & reg386[(4'hb):(4'hb)]) & (7'h41)) - $unsigned(forvar384));
            end
          reg396 <= $unsigned($unsigned((~|($unsigned(reg383) ?
              (^reg387) : reg386))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar397 = (1'h0); (forvar397 < (2'h3)); forvar397 = (forvar397 + (1'h1)))
        begin
          for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
            begin
              reg399 <= $signed(forvar384);
              reg400 = ({$signed((((8'hbd) ? reg392 : (8'ha3)) ?
                          ((8'hac) ? reg399 : reg393) : $unsigned(reg390)))} ?
                  ((!$signed(reg386[(1'h0):(1'h0)])) >> $signed((8'ha2))) : "Axo6ECcHHtnmO5zY8Lmw");
              reg401 <= $signed(forvar398);
              reg402 <= (8'hb7);
              reg403 <= ($unsigned((8'hb2)) ? "hWxXkxbDEoNk0y6" : wire375);
            end
          for (forvar404 = (1'h0); (forvar404 < (2'h2)); forvar404 = (forvar404 + (1'h1)))
            begin
              reg405 <= ($unsigned(wire375) ?
                  (reg386 << (reg387[(4'he):(4'hb)] ?
                      reg399 : (&wire377[(4'hc):(1'h1)]))) : (wire375[(4'h8):(2'h3)] ?
                      $unsigned($signed($unsigned(wire376))) : (~&"IYWULkZ")));
              reg406 = $unsigned(({$unsigned(forvar384[(3'h4):(1'h1)])} | forvar381[(2'h3):(1'h1)]));
            end
        end
      reg407 <= (~^($unsigned($unsigned($signed(reg382))) == reg403[(1'h0):(1'h0)]));
      for (forvar408 = (1'h0); (forvar408 < (2'h2)); forvar408 = (forvar408 + (1'h1)))
        begin
          reg409 = reg390;
          reg410 <= ((wire375 >>> reg387) ?
              ((^~($unsigned(reg405) >> (reg402 ?
                  (8'ha4) : wire374))) != ("RX3Pp6XHad" ?
                  ("YOQgZCeJ9LB" ?
                      $signed((8'hbd)) : wire377) : (^reg390))) : $unsigned(("AXNBUt8CHxlHl3" || $unsigned({forvar398}))));
          reg411 <= wire379;
          for (forvar412 = (1'h0); (forvar412 < (2'h2)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 = (&reg393);
              reg414 = ((~^$unsigned($signed({reg406}))) << (wire375 ?
                  {$signed(reg391)} : {$unsigned("DIer")}));
            end
        end
      for (forvar415 = (1'h0); (forvar415 < (1'h1)); forvar415 = (forvar415 + (1'h1)))
        begin
          reg416 <= ((~^reg387[(1'h1):(1'h0)]) ?
              {((~^(forvar384 < reg388)) ?
                      reg392 : reg390[(3'h7):(2'h3)])} : $signed(wire378));
          reg417 <= reg385[(2'h3):(2'h3)];
          for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
            begin
              reg419 = ((reg411[(1'h0):(1'h0)] ?
                  {(wire379 ? $signed(reg400) : $signed((8'hbe))),
                      $signed($unsigned(reg413))} : $signed($unsigned(reg391))) & {$signed($signed($signed((8'hb2))))});
            end
          if (forvar398[(4'h8):(1'h1)])
            begin
              reg420 = reg414;
              reg421 <= $unsigned($signed(({(wire379 != reg400),
                      "3GtX3T5tdL9fK"} ?
                  "exHxpyiKTqOflSutX4Qi" : {(reg387 ? forvar415 : wire379),
                      wire375[(4'hd):(3'h5)]})));
              reg422 <= {$signed(reg400)};
              reg423 <= $unsigned($signed("Rg5egP"));
            end
          else
            begin
              reg420 <= ({$signed(({reg391, reg387} || $unsigned(reg417))),
                  ((reg417 ?
                      (forvar397 - (7'h43)) : $unsigned(reg410)) ^~ $signed($signed(reg420)))} >> (forvar397[(2'h3):(2'h3)] <<< (!reg420)));
              reg421 = $unsigned($unsigned(forvar404));
            end
        end
    end
  always
    @(posedge clk) begin
      reg424 <= reg406;
      reg425 <= {(reg422[(2'h2):(2'h2)] ^ reg392[(5'h10):(1'h1)])};
      for (forvar426 = (1'h0); (forvar426 < (3'h4)); forvar426 = (forvar426 + (1'h1)))
        begin
          for (forvar427 = (1'h0); (forvar427 < (1'h0)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= (-(reg419[(3'h7):(1'h1)] >= reg393[(2'h2):(1'h1)]));
              reg429 = $signed({$unsigned((~^reg395[(3'h4):(1'h1)]))});
              reg430 <= ({forvar397} * (reg423[(4'hd):(3'h7)] ?
                  reg405[(2'h2):(1'h1)] : $unsigned("uWoKt9")));
              reg431 = $signed($unsigned(forvar384));
              reg432 = (8'hbe);
            end
        end
      if ($unsigned("TrRfdAF2NOEwk"))
        begin
          if ((reg394[(2'h2):(1'h1)] ?
              $signed((+(^~(forvar427 ?
                  reg410 : reg406)))) : (forvar412 & (&(reg417[(2'h2):(1'h0)] + (wire379 ?
                  reg416 : reg421))))))
            begin
              reg433 = $unsigned(forvar397[(2'h3):(1'h1)]);
            end
          else
            begin
              reg433 = (^$signed(forvar398[(2'h2):(1'h1)]));
              reg434 = (wire376 ?
                  $signed(reg400) : ($unsigned(((-reg414) ?
                          forvar397[(2'h3):(1'h0)] : (8'h9e))) ?
                      ((!$signed((7'h44))) > (reg388 <= reg399[(4'hc):(2'h2)])) : {($unsigned(reg399) >>> (~^reg385)),
                          $signed((-forvar426))}));
            end
          reg435 <= ((!$signed(reg410)) ?
              $unsigned({{reg409}, $signed(reg434)}) : ((reg432[(4'hd):(3'h6)] ?
                  reg380[(3'h6):(3'h6)] : reg386) && ($signed((reg410 ?
                      reg419 : (8'hb6))) ?
                  {(forvar398 >= wire375), reg387} : ((reg405 ?
                      (7'h44) : forvar398) != reg428))));
        end
      else
        begin
          for (forvar433 = (1'h0); (forvar433 < (1'h1)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= reg390[(2'h3):(1'h0)];
              reg435 <= reg388[(2'h3):(1'h0)];
            end
          for (forvar436 = (1'h0); (forvar436 < (1'h1)); forvar436 = (forvar436 + (1'h1)))
            begin
              reg437 = $signed(reg421[(4'he):(1'h1)]);
            end
          reg438 <= (((((~&reg413) <<< (~&(8'hb1))) ?
              (reg400[(2'h3):(1'h1)] && (reg420 - reg428)) : $signed((&reg413))) << (~((reg414 * reg406) ?
              (reg402 >= forvar426) : $signed(wire379)))) ~^ (!(&forvar426)));
          for (forvar439 = (1'h0); (forvar439 < (1'h1)); forvar439 = (forvar439 + (1'h1)))
            begin
              reg440 = $unsigned({(($unsigned(reg385) ?
                      forvar381[(4'hc):(4'hb)] : $unsigned(wire376)) - $signed(((8'hae) & reg396))),
                  $unsigned($unsigned(reg389[(1'h1):(1'h1)]))});
              reg441 = ((+"") ?
                  ({$signed($signed(reg425)),
                          {reg405[(2'h3):(1'h0)], {(8'ha6)}}} ?
                      reg411[(3'h5):(1'h0)] : $unsigned(({reg424} ?
                          reg423 : {(8'hb2),
                              forvar426}))) : reg410[(3'h4):(3'h4)]);
              reg442 <= ({($signed(reg417) ?
                      ((reg396 * reg406) ?
                          reg390[(1'h1):(1'h0)] : forvar412[(1'h1):(1'h1)]) : $signed($signed(reg387))),
                  reg382} >> {((8'ha2) ?
                      $signed((|reg422)) : reg402[(4'h9):(1'h0)]),
                  forvar415[(3'h5):(1'h1)]});
            end
        end
    end
  assign wire443 = {(~|"HyMNlLgaEMZP2Y3v9Q"), reg440};
  always
    @(posedge clk) begin
      for (forvar444 = (1'h0); (forvar444 < (1'h0)); forvar444 = (forvar444 + (1'h1)))
        begin
          for (forvar445 = (1'h0); (forvar445 < (1'h1)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= $unsigned(((~reg402[(4'hc):(2'h2)]) ?
                  $signed((-(reg410 && reg382))) : (8'h9d)));
              reg447 = $unsigned(forvar436[(2'h2):(1'h1)]);
            end
          for (forvar448 = (1'h0); (forvar448 < (1'h1)); forvar448 = (forvar448 + (1'h1)))
            begin
              reg449 = reg385[(2'h3):(1'h0)];
              reg450 = ((~&(-reg434[(2'h3):(1'h0)])) < {"Rfx7RQDbn6RlKnIOa"});
              reg451 = forvar408[(2'h3):(2'h2)];
              reg452 = (forvar426[(1'h1):(1'h1)] ?
                  (reg401 ?
                      reg403[(1'h1):(1'h1)] : $signed(reg402[(3'h4):(1'h1)])) : (reg392[(2'h2):(1'h0)] | forvar418));
              reg453 <= (~$unsigned($unsigned(($unsigned(reg428) + reg401))));
            end
          if ($signed($signed($signed((forvar439[(2'h2):(1'h0)] ?
              $signed(reg434) : (reg402 || forvar397))))))
            begin
              reg454 = ((wire443[(2'h3):(2'h2)] ?
                  ((~|reg401[(4'h9):(4'h8)]) ?
                      {$unsigned(reg387),
                          (reg393 ?
                              reg451 : reg453)} : reg449) : $unsigned($unsigned(reg416))) ~^ reg453);
              reg455 <= (reg416[(2'h3):(1'h0)] ?
                  {(wire374 ?
                          $unsigned((forvar404 * reg433)) : reg434[(3'h7):(2'h3)]),
                      $signed(reg405[(1'h0):(1'h0)])} : ((-{(~reg440)}) ?
                      (^$unsigned($unsigned(reg453))) : ({reg399} && (8'ha8))));
              reg456 <= $signed(reg416[(2'h3):(2'h2)]);
              reg457 <= ($signed($signed($signed((reg421 == (8'hbb))))) ?
                  (7'h44) : $unsigned($signed(($unsigned((8'ha1)) ?
                      (reg414 ? reg399 : reg456) : $unsigned(forvar404)))));
            end
          else
            begin
              reg454 <= $signed(((~reg425) ?
                  (reg438 != reg383[(2'h2):(1'h0)]) : reg399[(4'hc):(3'h6)]));
              reg455 <= ({reg442} ?
                  reg406[(4'ha):(2'h2)] : reg393[(1'h1):(1'h0)]);
            end
          reg458 <= (~|((-(+(reg442 ?
              reg417 : reg433))) > $unsigned(((reg440 ~^ wire374) >>> forvar427[(4'hd):(4'h8)]))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module173  (y, clk, wire178, wire177, wire176, wire175, wire174);
  output wire [(32'h8ec):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire178;
  input wire [(5'h14):(1'h0)] wire177;
  input wire [(5'h11):(1'h0)] wire176;
  input wire signed [(3'h4):(1'h0)] wire175;
  input wire [(4'hc):(1'h0)] wire174;
  wire [(2'h2):(1'h0)] wire370;
  wire [(5'h11):(1'h0)] wire369;
  wire signed [(3'h7):(1'h0)] wire368;
  wire [(4'hc):(1'h0)] wire367;
  wire [(4'h9):(1'h0)] wire366;
  wire signed [(3'h4):(1'h0)] wire365;
  wire [(3'h6):(1'h0)] wire364;
  reg signed [(4'hd):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg362 = (1'h0);
  reg [(4'ha):(1'h0)] reg361 = (1'h0);
  reg [(4'hc):(1'h0)] reg360 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg359 = (1'h0);
  reg [(4'hd):(1'h0)] reg358 = (1'h0);
  reg [(4'ha):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar356 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg355 = (1'h0);
  reg [(3'h4):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg352 = (1'h0);
  reg [(5'h11):(1'h0)] forvar351 = (1'h0);
  reg [(4'hf):(1'h0)] reg350 = (1'h0);
  reg [(4'hb):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg348 = (1'h0);
  reg [(5'h11):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg345 = (1'h0);
  reg [(5'h12):(1'h0)] reg344 = (1'h0);
  reg [(5'h13):(1'h0)] reg343 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg342 = (1'h0);
  reg [(4'hd):(1'h0)] forvar341 = (1'h0);
  reg [(3'h4):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg339 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg338 = (1'h0);
  reg [(4'he):(1'h0)] forvar337 = (1'h0);
  reg [(5'h12):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg335 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar334 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar333 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire332;
  reg [(2'h2):(1'h0)] reg331 = (1'h0);
  reg [(5'h13):(1'h0)] reg330 = (1'h0);
  reg [(4'h9):(1'h0)] reg329 = (1'h0);
  reg [(5'h12):(1'h0)] reg328 = (1'h0);
  reg [(4'h8):(1'h0)] reg327 = (1'h0);
  reg [(4'hd):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar325 = (1'h0);
  reg [(4'h8):(1'h0)] reg324 = (1'h0);
  reg [(4'hf):(1'h0)] reg323 = (1'h0);
  reg [(4'hf):(1'h0)] reg322 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg321 = (1'h0);
  reg [(2'h2):(1'h0)] reg320 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar319 = (1'h0);
  reg [(2'h3):(1'h0)] reg318 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg317 = (1'h0);
  reg [(4'ha):(1'h0)] reg316 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar314 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg312 = (1'h0);
  reg [(4'hc):(1'h0)] reg311 = (1'h0);
  reg [(5'h11):(1'h0)] reg310 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg308 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg306 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg305 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar304 = (1'h0);
  reg [(4'h8):(1'h0)] reg303 = (1'h0);
  reg [(3'h5):(1'h0)] reg302 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar301 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar300 = (1'h0);
  wire [(3'h6):(1'h0)] wire299;
  wire signed [(3'h6):(1'h0)] wire298;
  reg [(4'hb):(1'h0)] reg297 = (1'h0);
  reg [(5'h11):(1'h0)] reg296 = (1'h0);
  reg [(4'h8):(1'h0)] forvar295 = (1'h0);
  reg [(3'h5):(1'h0)] reg294 = (1'h0);
  reg [(2'h3):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg291 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg290 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg288 = (1'h0);
  reg [(5'h11):(1'h0)] reg287 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar285 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar284 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg283 = (1'h0);
  reg [(4'h9):(1'h0)] reg282 = (1'h0);
  reg [(5'h12):(1'h0)] reg281 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg280 = (1'h0);
  reg [(5'h10):(1'h0)] reg279 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar278 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg277 = (1'h0);
  reg [(5'h12):(1'h0)] forvar276 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg275 = (1'h0);
  reg [(2'h3):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar270 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg269 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg267 = (1'h0);
  reg [(4'h8):(1'h0)] reg266 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg265 = (1'h0);
  reg [(2'h3):(1'h0)] reg264 = (1'h0);
  reg [(5'h15):(1'h0)] forvar263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar260 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg259 = (1'h0);
  reg [(4'hf):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(5'h12):(1'h0)] reg256 = (1'h0);
  reg [(4'he):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar254 = (1'h0);
  reg [(3'h4):(1'h0)] reg253 = (1'h0);
  reg [(5'h15):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg249 = (1'h0);
  reg [(5'h10):(1'h0)] forvar248 = (1'h0);
  reg [(4'hd):(1'h0)] forvar247 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg246 = (1'h0);
  reg [(4'hc):(1'h0)] forvar245 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg242 = (1'h0);
  reg [(4'hb):(1'h0)] forvar241 = (1'h0);
  reg [(4'hf):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg238 = (1'h0);
  reg [(5'h15):(1'h0)] reg237 = (1'h0);
  reg [(4'he):(1'h0)] forvar236 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar235 = (1'h0);
  reg [(4'h9):(1'h0)] reg234 = (1'h0);
  reg [(4'h8):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg232 = (1'h0);
  reg [(4'h9):(1'h0)] reg231 = (1'h0);
  reg [(5'h11):(1'h0)] reg230 = (1'h0);
  reg [(4'hd):(1'h0)] forvar229 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar228 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg227 = (1'h0);
  reg [(5'h10):(1'h0)] reg226 = (1'h0);
  reg [(2'h3):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar222 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg218 = (1'h0);
  reg [(5'h10):(1'h0)] reg217 = (1'h0);
  reg [(4'ha):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg215 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar213 = (1'h0);
  reg [(4'hc):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg211 = (1'h0);
  reg [(4'h8):(1'h0)] reg210 = (1'h0);
  reg [(3'h7):(1'h0)] reg209 = (1'h0);
  reg [(3'h7):(1'h0)] forvar208 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar207 = (1'h0);
  reg [(4'hb):(1'h0)] reg206 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg205 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg204 = (1'h0);
  reg [(4'hf):(1'h0)] reg203 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg202 = (1'h0);
  reg [(4'hb):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg199 = (1'h0);
  reg [(3'h5):(1'h0)] reg198 = (1'h0);
  reg [(5'h14):(1'h0)] reg197 = (1'h0);
  reg [(2'h3):(1'h0)] forvar196 = (1'h0);
  reg [(4'hd):(1'h0)] reg195 = (1'h0);
  reg [(3'h6):(1'h0)] forvar194 = (1'h0);
  wire [(4'ha):(1'h0)] wire193;
  wire [(4'hf):(1'h0)] wire192;
  wire [(5'h12):(1'h0)] wire191;
  reg [(3'h7):(1'h0)] reg190 = (1'h0);
  reg [(4'ha):(1'h0)] reg189 = (1'h0);
  reg [(5'h13):(1'h0)] reg188 = (1'h0);
  reg [(4'he):(1'h0)] reg187 = (1'h0);
  reg [(5'h13):(1'h0)] forvar186 = (1'h0);
  reg [(5'h15):(1'h0)] reg184 = (1'h0);
  reg [(4'hf):(1'h0)] forvar182 = (1'h0);
  reg [(3'h6):(1'h0)] reg185 = (1'h0);
  reg [(4'ha):(1'h0)] forvar184 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg183 = (1'h0);
  reg [(4'h9):(1'h0)] reg182 = (1'h0);
  reg [(4'hf):(1'h0)] reg181 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire180;
  wire signed [(3'h7):(1'h0)] wire179;
  assign y = {wire370,
                 wire369,
                 wire368,
                 wire367,
                 wire366,
                 wire365,
                 wire364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 forvar356,
                 reg355,
                 reg351,
                 reg354,
                 reg353,
                 reg352,
                 forvar351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 forvar346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 forvar341,
                 reg340,
                 reg339,
                 reg338,
                 forvar337,
                 reg336,
                 reg335,
                 forvar334,
                 forvar333,
                 wire332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 forvar325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 forvar319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 forvar314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 forvar309,
                 reg308,
                 forvar307,
                 reg306,
                 reg305,
                 forvar304,
                 reg303,
                 reg302,
                 forvar301,
                 forvar300,
                 wire299,
                 wire298,
                 reg297,
                 reg296,
                 forvar295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 forvar285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 forvar278,
                 reg277,
                 forvar276,
                 reg275,
                 reg263,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 reg261,
                 forvar260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 forvar254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 forvar248,
                 forvar247,
                 reg246,
                 forvar245,
                 reg244,
                 reg243,
                 reg242,
                 forvar241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 forvar236,
                 forvar235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 forvar229,
                 forvar228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 forvar222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 forvar213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 forvar208,
                 forvar207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 forvar196,
                 reg195,
                 forvar194,
                 wire193,
                 wire192,
                 wire191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 forvar186,
                 reg184,
                 forvar182,
                 reg185,
                 forvar184,
                 reg183,
                 reg182,
                 reg181,
                 wire180,
                 wire179,
                 (1'h0)};
  assign wire179 = $signed(wire176[(1'h0):(1'h0)]);
  assign wire180 = ($unsigned($signed({(~^wire176),
                       (8'hb5)})) - ($signed($signed((wire179 ?
                           (7'h40) : wire178))) ?
                       $unsigned($signed($signed((8'hbb)))) : {wire175,
                           (((7'h40) != wire178) <= wire179)}));
  always
    @(posedge clk) begin
      if ($signed((|(wire175[(3'h4):(2'h2)] == {wire180,
          (wire178 ? wire177 : wire178)}))))
        begin
          if ((|$unsigned(wire180[(1'h0):(1'h0)])))
            begin
              reg181 <= ({$unsigned(wire180[(2'h3):(1'h1)])} > $signed($signed(($signed(wire175) ?
                  $signed(wire175) : wire176[(3'h6):(1'h0)]))));
              reg182 <= wire179[(2'h2):(1'h0)];
              reg183 = (^~(wire175[(1'h1):(1'h0)] + $unsigned("xhLbWPBTsra8TwLSGah")));
            end
          else
            begin
              reg181 <= reg183[(1'h0):(1'h0)];
              reg182 = "eqUF";
            end
          for (forvar184 = (1'h0); (forvar184 < (2'h2)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 <= ((~^({wire177} & (&$signed(reg181)))) ?
                  "2g76kzGYbhFv" : {$signed($unsigned((8'hbc))),
                      wire178[(3'h4):(3'h4)]});
            end
        end
      else
        begin
          reg181 = ((wire180 >> (((wire177 ?
              wire176 : wire176) >>> $signed(reg181)) & ($unsigned(reg181) ?
              (~reg181) : reg183))) < (~&{($signed(wire179) ?
                  (reg183 ? wire177 : forvar184) : (+reg181)),
              wire179}));
          for (forvar182 = (1'h0); (forvar182 < (1'h0)); forvar182 = (forvar182 + (1'h1)))
            begin
              reg183 <= wire179;
              reg184 = ((8'ha2) ? forvar182 : ($unsigned(wire174) ^ reg185));
              reg185 = (&($unsigned($signed((wire179 ? reg184 : reg181))) ?
                  (~^$unsigned($signed(wire175))) : $signed($signed(wire179[(2'h3):(1'h0)]))));
            end
          for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg187 = ((|$signed(((|reg182) ?
                      $signed((8'h9d)) : (&wire174)))) ?
                  forvar184[(3'h7):(2'h2)] : wire177);
              reg188 = wire177;
              reg189 <= (|reg182);
              reg190 = ($signed($signed(wire175[(2'h2):(2'h2)])) ?
                  (~^$signed((wire180 ?
                      $signed(reg185) : (forvar184 >> forvar184)))) : {(-((8'ha8) ~^ (~forvar184)))});
            end
        end
    end
  assign wire191 = {$signed(reg189)};
  assign wire192 = wire178;
  assign wire193 = reg187[(4'h9):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar194 = (1'h0); (forvar194 < (1'h0)); forvar194 = (forvar194 + (1'h1)))
        begin
          reg195 = $signed($unsigned((("memPYXAnOcvA0HKWRPgh" ?
              (reg188 ?
                  reg183 : (8'h9f)) : $unsigned(reg182)) || $signed(reg188[(4'h9):(2'h2)]))));
          for (forvar196 = (1'h0); (forvar196 < (1'h1)); forvar196 = (forvar196 + (1'h1)))
            begin
              reg197 = forvar184[(3'h4):(1'h0)];
              reg198 = wire191;
              reg199 <= $signed((~&{((forvar194 ? wire192 : wire193) ~^ reg190),
                  $unsigned(reg184)}));
              reg200 <= (&(~^{forvar182, $unsigned($unsigned(wire174))}));
            end
          reg201 = (!$signed({((reg185 ? reg200 : wire191) ?
                  (wire175 ? forvar194 : reg200) : (reg197 ?
                      wire180 : forvar186)),
              reg195}));
          reg202 = $signed((((&$unsigned((8'hbd))) ?
                  $signed((wire174 ?
                      reg182 : wire175)) : reg181[(2'h3):(1'h1)]) ?
              reg195[(4'h9):(3'h6)] : reg189));
          if ((((~&$signed(forvar196[(2'h3):(1'h0)])) ?
                  $signed(reg195[(3'h7):(3'h6)]) : "59puh0s9TPZNbN32zgk6") ?
              {forvar196[(2'h3):(1'h1)]} : ((wire192[(2'h3):(2'h2)] ?
                  {(reg181 >>> reg183)} : $unsigned(wire180)) ~^ wire193)))
            begin
              reg203 = $unsigned($signed((~&forvar182[(4'hf):(1'h1)])));
            end
          else
            begin
              reg203 = (^~($unsigned(($unsigned(forvar186) - {reg184,
                      reg187})) ?
                  wire178 : reg202));
              reg204 <= (~{(wire177 ^ reg183), forvar196[(2'h2):(1'h1)]});
              reg205 <= reg203[(4'hf):(1'h1)];
              reg206 = $unsigned($unsigned({""}));
            end
        end
      for (forvar207 = (1'h0); (forvar207 < (2'h2)); forvar207 = (forvar207 + (1'h1)))
        begin
          for (forvar208 = (1'h0); (forvar208 < (2'h3)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 <= (wire192 ?
                  (wire178 ?
                      ({$unsigned((8'hbc))} >= (((8'ha5) && wire179) >= $signed(wire178))) : $unsigned(forvar184)) : wire177[(1'h1):(1'h0)]);
              reg210 <= (((reg200 ?
                          (reg201 | (wire180 ?
                              reg190 : reg181)) : ($signed(reg182) ?
                              (~forvar182) : reg202)) ?
                      reg204 : ($signed(reg206) >> ($unsigned(reg205) ?
                          wire177[(4'hb):(4'h9)] : $signed((8'hb9))))) ?
                  "" : wire178);
              reg211 <= ($signed($signed(forvar182[(3'h4):(2'h3)])) * $signed({(+$signed((7'h41)))}));
              reg212 = (({(reg190[(3'h4):(3'h4)] * (+reg203)),
                  $signed({reg202})} ^ ({$signed(reg189)} * $unsigned({wire193,
                  forvar196}))) <<< $signed(forvar196));
            end
          for (forvar213 = (1'h0); (forvar213 < (1'h0)); forvar213 = (forvar213 + (1'h1)))
            begin
              reg214 = forvar194;
              reg215 = ($signed(reg211) ?
                  wire177[(4'h8):(2'h2)] : {(-(reg188[(3'h7):(1'h1)] >> (-wire175)))});
            end
          reg216 = reg200;
          if ({$signed($unsigned(reg185)),
              ($signed(reg204) ?
                  $signed($signed($unsigned(wire177))) : wire179)})
            begin
              reg217 <= reg202;
              reg218 <= ({(-((8'hbc) ?
                      (reg204 | reg216) : (~^wire180)))} >> ($signed((-(!(8'ha7)))) <<< $signed($unsigned(reg210[(2'h3):(1'h1)]))));
              reg219 = (wire176 <<< (reg198 < "XIgoKe2sB"));
              reg220 = (|{($unsigned((wire191 || reg200)) ?
                      "yce610CDGw" : ((reg205 || reg203) && $signed(reg202))),
                  reg185[(1'h1):(1'h0)]});
              reg221 <= reg198;
            end
          else
            begin
              reg217 = $unsigned((8'hbd));
              reg218 <= wire191[(2'h3):(2'h3)];
            end
          for (forvar222 = (1'h0); (forvar222 < (2'h3)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 = reg214[(1'h1):(1'h0)];
              reg224 <= (~$unsigned((&$unsigned(reg212))));
              reg225 <= (~&($unsigned((~|(wire179 < reg197))) <<< (-reg212)));
              reg226 = {("I0Xr" ?
                      $unsigned(($signed(wire180) ?
                          wire179[(3'h4):(2'h2)] : {(8'hbc),
                              reg219})) : wire177[(5'h11):(4'he)]),
                  $unsigned(reg198[(2'h3):(2'h2)])};
              reg227 = $unsigned({((^~(reg201 ?
                      reg197 : wire175)) != $unsigned(forvar184[(1'h0):(1'h0)]))});
            end
        end
      for (forvar228 = (1'h0); (forvar228 < (2'h2)); forvar228 = (forvar228 + (1'h1)))
        begin
          for (forvar229 = (1'h0); (forvar229 < (3'h4)); forvar229 = (forvar229 + (1'h1)))
            begin
              reg230 <= reg198[(3'h5):(3'h4)];
              reg231 <= {$signed({(~reg195),
                      (reg230[(4'ha):(3'h7)] ?
                          {wire192, reg206} : reg223[(1'h0):(1'h0)])})};
              reg232 <= ($unsigned(((~^((8'hb5) << wire180)) ~^ ($unsigned(reg211) ?
                  (7'h41) : $unsigned(wire177)))) || $unsigned((((+forvar196) + (reg187 * wire176)) << "32ygG1x1N6ACmBkAY")));
              reg233 = (+$signed((($signed(reg202) ?
                  $signed(reg211) : reg199[(4'h8):(3'h5)]) || $signed($unsigned(reg223)))));
              reg234 <= ($signed(reg232[(4'h8):(1'h0)]) <<< reg233);
            end
        end
      for (forvar235 = (1'h0); (forvar235 < (2'h3)); forvar235 = (forvar235 + (1'h1)))
        begin
          for (forvar236 = (1'h0); (forvar236 < (1'h1)); forvar236 = (forvar236 + (1'h1)))
            begin
              reg237 <= ((wire192 > {$signed(reg215[(1'h1):(1'h0)])}) ?
                  (wire174[(3'h7):(1'h1)] - reg220[(3'h4):(2'h2)]) : reg214[(1'h0):(1'h0)]);
              reg238 <= ({$signed(($signed(reg227) * (|reg197)))} && $signed(forvar208));
              reg239 <= ((!(~|((reg220 == wire191) ?
                  reg237 : (~|reg181)))) > ((reg185[(1'h0):(1'h0)] == $unsigned(reg216[(4'ha):(2'h3)])) ?
                  reg218[(2'h3):(2'h2)] : reg211[(4'he):(4'h8)]));
              reg240 = reg185;
            end
          for (forvar241 = (1'h0); (forvar241 < (3'h4)); forvar241 = (forvar241 + (1'h1)))
            begin
              reg242 <= $unsigned(wire175);
              reg243 <= (($signed(forvar228) || forvar208[(1'h0):(1'h0)]) ?
                  $unsigned($unsigned(((-reg219) ?
                      $signed(reg215) : reg227[(3'h6):(3'h4)]))) : (~(8'hab)));
            end
          reg244 = (~&reg214);
          for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
            begin
              reg246 <= reg210;
            end
        end
      for (forvar247 = (1'h0); (forvar247 < (3'h4)); forvar247 = (forvar247 + (1'h1)))
        begin
          for (forvar248 = (1'h0); (forvar248 < (1'h1)); forvar248 = (forvar248 + (1'h1)))
            begin
              reg249 <= {((8'ha9) ?
                      $unsigned((+(forvar184 ?
                          reg243 : wire178))) : ((7'h44) == wire176)),
                  $signed($signed((forvar228 ?
                      $unsigned(wire177) : (reg187 && (8'hb4)))))};
              reg250 <= ($unsigned($signed(({wire180} ?
                      $signed((7'h44)) : $unsigned(reg233)))) ?
                  "k2p7RZZkwbHrEoDk" : ((forvar194 ?
                      "PCtlu23m2PM" : $signed({reg189})) ^ $unsigned(({wire176} ?
                      reg205[(1'h0):(1'h0)] : (forvar194 ? reg212 : reg198)))));
              reg251 <= reg201;
              reg252 = ($signed($signed($unsigned(wire192[(2'h3):(1'h0)]))) < (~^reg185[(3'h6):(3'h4)]));
              reg253 <= $unsigned(((({forvar241} ?
                  (reg189 << wire175) : $signed(reg238)) ~^ ((reg211 != reg231) ?
                  reg252 : (reg189 ?
                      reg209 : reg200))) | "liizEnZhMo5QmIsk1TYw"));
            end
          for (forvar254 = (1'h0); (forvar254 < (2'h3)); forvar254 = (forvar254 + (1'h1)))
            begin
              reg255 <= wire176;
              reg256 = $unsigned(forvar235[(3'h4):(3'h4)]);
              reg257 = ($signed(wire178[(3'h4):(1'h0)]) | forvar213[(1'h0):(1'h0)]);
              reg258 = (forvar182[(3'h7):(1'h1)] ?
                  (reg230[(4'ha):(3'h4)] ?
                      wire193[(3'h7):(3'h5)] : reg219[(1'h1):(1'h0)]) : reg181[(1'h1):(1'h0)]);
            end
          reg259 <= reg206;
          for (forvar260 = (1'h0); (forvar260 < (2'h3)); forvar260 = (forvar260 + (1'h1)))
            begin
              reg261 = $unsigned((^({reg206[(2'h3):(2'h3)]} ?
                  $signed({reg239, forvar248}) : ("CpBFF2Aaicg5XHId" ?
                      $signed(wire175) : reg243))));
              reg262 = (~|(^{reg203, (8'ha4)}));
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg201[(2'h3):(1'h1)])
        begin
          for (forvar263 = (1'h0); (forvar263 < (2'h2)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 <= ($signed((8'hb6)) ?
                  $unsigned((forvar213[(2'h2):(2'h2)] <<< ($signed(reg204) ?
                      reg182[(3'h4):(1'h0)] : (reg214 * forvar254)))) : $unsigned(($signed(((8'hbb) ?
                          (8'ha5) : reg182)) ?
                      (8'ha1) : ({reg187} ? (-reg197) : (reg233 * reg224)))));
              reg265 = reg181[(2'h2):(1'h1)];
              reg266 <= {(reg253 ?
                      reg227[(2'h2):(2'h2)] : $signed((reg182[(3'h4):(1'h1)] ?
                          reg212[(2'h2):(2'h2)] : (^reg211)))),
                  (((forvar207 && $signed(reg231)) << reg216) ?
                      reg211 : $signed({(reg238 ^ forvar229), (|reg201)}))};
              reg267 <= $signed(reg244[(3'h6):(3'h4)]);
              reg268 = $signed({$unsigned($unsigned((^wire174)))});
            end
          reg269 = ((((wire192 ? $signed(reg183) : $signed(reg195)) - reg188) ?
              (8'hba) : $signed((~|((8'ha2) * reg230)))) ^~ (!$signed(reg182[(2'h2):(1'h1)])));
          for (forvar270 = (1'h0); (forvar270 < (2'h2)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 = reg261[(2'h2):(1'h1)];
              reg272 <= (($unsigned(reg257) ?
                      (($unsigned(wire174) & $signed((7'h44))) & reg200) : reg199) ?
                  reg261[(2'h2):(1'h0)] : $unsigned($signed((^~$unsigned(reg239)))));
              reg273 = (reg224 <= {($unsigned(reg255) ?
                      $signed((-reg237)) : ""),
                  {($signed(reg230) ? reg184 : {(8'hb8), reg251})}});
            end
          reg274 <= (&{($signed((reg223 * reg257)) - $unsigned($signed(reg255)))});
        end
      else
        begin
          if (reg268[(1'h1):(1'h0)])
            begin
              reg263 = ($unsigned((~^$signed(reg198[(3'h4):(3'h4)]))) ?
                  (~|($signed($unsigned((8'haa))) > $unsigned(reg218[(3'h6):(3'h5)]))) : (+("VUus" ^ (reg251[(4'h9):(3'h5)] ?
                      $unsigned(reg185) : forvar229))));
              reg264 = $signed(((~($signed(reg205) ?
                      (reg212 ? reg264 : (8'haf)) : (reg271 ?
                          wire193 : forvar235))) ?
                  $unsigned((~&reg274[(3'h4):(1'h0)])) : $unsigned($unsigned($signed((8'ha1))))));
            end
          else
            begin
              reg263 = (reg243 ? reg264[(1'h0):(1'h0)] : (7'h40));
            end
        end
      reg275 = $unsigned((!wire175[(1'h1):(1'h1)]));
      for (forvar276 = (1'h0); (forvar276 < (3'h4)); forvar276 = (forvar276 + (1'h1)))
        begin
          reg277 = reg181;
          for (forvar278 = (1'h0); (forvar278 < (2'h2)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 = $unsigned({$signed(((reg205 ?
                      reg187 : forvar194) * $signed(reg215)))});
              reg280 <= ((~$signed(reg209[(1'h0):(1'h0)])) ? reg231 : reg249);
              reg281 <= (8'hae);
            end
          reg282 <= {$signed(reg256)};
          reg283 = ($unsigned(forvar260[(2'h2):(2'h2)]) >> {reg263});
        end
      for (forvar284 = (1'h0); (forvar284 < (1'h1)); forvar284 = (forvar284 + (1'h1)))
        begin
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 <= reg250;
              reg287 = reg252[(4'ha):(1'h1)];
              reg288 = reg211;
            end
          reg289 <= reg209[(3'h5):(2'h3)];
          reg290 = ($signed({$unsigned($unsigned(reg221)),
                  ($unsigned((8'haa)) ? (^reg283) : (reg238 <= wire176))}) ?
              $unsigned((reg243 ?
                  forvar284[(4'he):(3'h7)] : reg206[(4'ha):(3'h7)])) : forvar254[(4'h8):(3'h5)]);
          if ((&forvar228))
            begin
              reg291 <= $signed((~^(^~forvar254)));
              reg292 <= reg203[(3'h6):(2'h2)];
              reg293 <= wire176[(4'hc):(3'h4)];
              reg294 <= $signed(((~|"aft1IC2") ?
                  reg249 : {$signed((reg233 ? wire177 : (8'ha1))),
                      (((8'hbe) ? reg211 : reg289) ?
                          reg240[(3'h7):(3'h6)] : (wire175 ?
                              (8'hab) : reg211))}));
            end
          else
            begin
              reg291 = $signed($signed($signed(((reg264 ? wire193 : reg219) ?
                  reg184 : (-reg252)))));
              reg292 = (&((8'hbb) ?
                  (forvar207 ?
                      $signed(reg231[(2'h3):(1'h1)]) : reg234) : ((~$signed(forvar208)) | forvar186[(4'hc):(3'h4)])));
              reg293 <= reg272[(4'hb):(2'h3)];
              reg294 <= (reg189[(4'h9):(4'h9)] << $unsigned($signed({reg275[(4'hc):(2'h3)],
                  reg289})));
            end
          for (forvar295 = (1'h0); (forvar295 < (2'h2)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 = reg251;
            end
        end
    end
  always
    @(posedge clk) begin
      reg297 = forvar184;
    end
  assign wire298 = (((((&(8'ha9)) ?
                           $signed(reg293) : $unsigned(reg215)) ~^ $signed(reg210)) - (reg206[(3'h5):(1'h0)] ?
                           {(reg275 ? reg266 : reg252),
                               $signed(forvar228)} : $signed($unsigned(reg291)))) ?
                       $signed(reg243) : reg292[(3'h5):(2'h3)]);
  assign wire299 = forvar229;
  always
    @(posedge clk) begin
      for (forvar300 = (1'h0); (forvar300 < (1'h1)); forvar300 = (forvar300 + (1'h1)))
        begin
          for (forvar301 = (1'h0); (forvar301 < (1'h1)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= forvar285;
              reg303 = $unsigned(reg288[(5'h14):(4'hc)]);
            end
          for (forvar304 = (1'h0); (forvar304 < (1'h0)); forvar304 = (forvar304 + (1'h1)))
            begin
              reg305 = reg280[(2'h3):(2'h3)];
            end
          reg306 = {$signed({((reg224 ? reg244 : forvar194) ?
                      $signed(forvar247) : {reg205, reg293}),
                  $signed(reg289)}),
              reg282};
        end
      for (forvar307 = (1'h0); (forvar307 < (2'h2)); forvar307 = (forvar307 + (1'h1)))
        begin
          reg308 = forvar241;
          for (forvar309 = (1'h0); (forvar309 < (3'h4)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 <= $unsigned(reg259);
              reg311 <= (7'h40);
              reg312 <= (8'ha5);
            end
          reg313 <= {$unsigned((^{reg226[(3'h7):(3'h6)],
                  (forvar241 ? reg210 : reg239)})),
              (wire191[(5'h11):(4'hc)] ?
                  $unsigned($signed(reg262)) : ($unsigned($signed(reg251)) ?
                      $signed(reg280[(1'h1):(1'h0)]) : $unsigned(reg306)))};
        end
      for (forvar314 = (1'h0); (forvar314 < (1'h1)); forvar314 = (forvar314 + (1'h1)))
        begin
          if (((!(forvar307 ?
              (+forvar229) : reg259)) ~^ ($unsigned($signed(reg246[(2'h2):(1'h0)])) ?
              $signed(reg250[(4'h9):(4'h8)]) : ($signed($signed(reg231)) && ((reg203 >> reg264) ?
                  $unsigned(wire178) : (+reg280))))))
            begin
              reg315 <= reg226[(4'hc):(2'h3)];
              reg316 <= {$signed($unsigned(reg237[(3'h7):(2'h3)])),
                  reg264[(2'h2):(1'h0)]};
            end
          else
            begin
              reg315 <= "q707X5vr5kwdDNG5gxq";
            end
          reg317 = {{$unsigned(reg240), $signed((~^(-reg316)))}};
          reg318 <= (($unsigned(((reg215 || forvar196) <<< wire179)) & {($unsigned((8'had)) ^~ (reg243 ?
                      reg261 : forvar208))}) ?
              ((($unsigned(forvar307) <= wire192[(1'h0):(1'h0)]) <= ((~^reg219) || $unsigned(forvar301))) >= (-((reg231 ^ forvar213) >>> wire180))) : (~(($signed(reg233) - $unsigned(reg292)) >= ("q1EBEDmLYB" ?
                  reg303 : (reg184 ? reg296 : (8'ha8))))));
        end
      for (forvar319 = (1'h0); (forvar319 < (2'h3)); forvar319 = (forvar319 + (1'h1)))
        begin
          reg320 <= $unsigned($unsigned($unsigned(((!forvar263) && $unsigned(reg230)))));
          if ($signed(reg282))
            begin
              reg321 = (8'ha1);
              reg322 <= $unsigned($unsigned((($signed((8'hb1)) >>> (|reg277)) ?
                  {(wire298 ? (8'hb9) : (8'hba))} : $unsigned(((8'hb2) ?
                      (8'hb0) : reg201)))));
              reg323 <= ((^~"THk") ^~ ($signed(wire177[(5'h10):(1'h0)]) ?
                  ($signed(forvar235[(3'h5):(1'h1)]) > (~^forvar254[(4'hf):(4'hd)])) : (|{$signed((8'hb6)),
                      (8'ha9)})));
            end
          else
            begin
              reg321 = reg201;
              reg322 <= $unsigned($signed($unsigned($signed(reg262[(3'h6):(3'h4)]))));
              reg323 <= (~^$signed(({(forvar182 & reg259),
                  $signed(reg302)} << (|forvar284))));
              reg324 <= ((!({"oDyPu"} ?
                      {reg257,
                          reg219[(1'h0):(1'h0)]} : (-(reg184 ~^ reg256)))) ?
                  {(($unsigned((7'h44)) << (forvar295 ^ forvar229)) ^ forvar247)} : $unsigned(reg318[(2'h2):(1'h1)]));
            end
          for (forvar325 = (1'h0); (forvar325 < (1'h0)); forvar325 = (forvar325 + (1'h1)))
            begin
              reg326 = (!{reg219[(2'h2):(1'h1)], {$unsigned(wire177)}});
            end
          if ((8'ha7))
            begin
              reg327 = {reg244[(5'h11):(1'h0)],
                  $unsigned({(+reg320), {(reg257 * (7'h42))}})};
              reg328 = reg209;
            end
          else
            begin
              reg327 <= (reg230[(3'h5):(2'h2)] ?
                  $unsigned(($signed(reg253) >> ((reg316 ?
                      reg230 : reg324) <<< (reg282 ?
                      reg282 : wire179)))) : $signed((({forvar186, wire298} ?
                      (~^reg262) : {reg240}) ^ (~|(reg282 << reg209)))));
              reg328 = $signed((~^$signed((~&(reg195 << (8'hb8))))));
              reg329 <= {$unsigned($signed((wire175 != {reg199, reg195}))),
                  (-(~|$unsigned((&(8'hbc)))))};
              reg330 <= {({(wire178[(3'h5):(3'h5)] ?
                          forvar184[(4'h8):(3'h5)] : {forvar194}),
                      $unsigned({reg292})} != reg198)};
            end
        end
      reg331 = ((~^((forvar186 && $unsigned((8'ha6))) ?
          ("YcH7v" ?
              $signed(wire174) : reg272[(5'h10):(4'hb)]) : $unsigned((reg243 ?
              (8'ha9) : forvar284)))) + $unsigned(reg261[(2'h2):(1'h1)]));
    end
  assign wire332 = ($signed((7'h41)) <= $unsigned($unsigned($unsigned($unsigned(reg197)))));
  always
    @(posedge clk) begin
      for (forvar333 = (1'h0); (forvar333 < (2'h3)); forvar333 = (forvar333 + (1'h1)))
        begin
          for (forvar334 = (1'h0); (forvar334 < (2'h2)); forvar334 = (forvar334 + (1'h1)))
            begin
              reg335 <= forvar245;
              reg336 = $unsigned(((((8'hb2) ?
                      {reg216,
                          reg280} : $unsigned(reg327)) ^ {(wire180 || forvar222)}) ?
                  (forvar285 ?
                      forvar248[(1'h1):(1'h0)] : $signed((-reg204))) : (8'ha5)));
            end
        end
      if (forvar325)
        begin
          for (forvar337 = (1'h0); (forvar337 < (3'h4)); forvar337 = (forvar337 + (1'h1)))
            begin
              reg338 = $unsigned((~^{{$signed(reg230)}}));
              reg339 <= $signed($signed(($unsigned(reg182[(2'h3):(1'h0)]) && reg282)));
              reg340 = $unsigned(("J" ?
                  (-($signed(reg246) > (8'had))) : (&(((8'h9f) ?
                          reg310 : reg279) ?
                      (forvar307 ?
                          (8'hb2) : reg286) : forvar270[(4'he):(3'h6)]))));
            end
          for (forvar341 = (1'h0); (forvar341 < (3'h4)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 <= $signed(((^~(&(7'h40))) ?
                  forvar301[(4'hd):(4'h9)] : reg219[(3'h4):(1'h0)]));
              reg343 = $unsigned((forvar304 ? reg275 : {$signed(forvar325)}));
              reg344 <= (8'ha9);
            end
          reg345 = "tVuOU5UqHEbTlBmw68CR";
          for (forvar346 = (1'h0); (forvar346 < (1'h0)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 = $unsigned(reg272[(2'h2):(1'h0)]);
              reg348 <= (-reg195);
              reg349 = $signed(forvar301);
            end
          reg350 = ($unsigned({reg264[(1'h0):(1'h0)],
              (+reg258[(4'ha):(1'h0)])}) != reg214);
        end
      else
        begin
          for (forvar337 = (1'h0); (forvar337 < (3'h4)); forvar337 = (forvar337 + (1'h1)))
            begin
              reg338 = reg231;
              reg339 = forvar284[(4'h8):(3'h7)];
            end
        end
      if (reg209)
        begin
          for (forvar351 = (1'h0); (forvar351 < (3'h4)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 = "VC3zShi";
              reg353 = $signed({(~|{$unsigned(reg203), (|reg210)})});
              reg354 = $signed((8'ha2));
            end
        end
      else
        begin
          if ((reg190[(3'h5):(3'h5)] ? reg233 : wire299[(3'h6):(2'h3)]))
            begin
              reg351 <= (reg224 ?
                  $unsigned((^({forvar284,
                      reg255} ^~ "JpzlKRv6MhZ"))) : reg353);
            end
          else
            begin
              reg351 <= (-$signed((forvar278[(4'hb):(1'h1)] << reg214)));
              reg352 <= "GIdv1R5Rny93fPn2lGK";
              reg353 <= (((wire176 ?
                      ((forvar351 * reg269) && (8'ha8)) : reg306) ?
                  $signed((reg321 || $unsigned(forvar208))) : {($signed(reg224) ?
                          (reg318 > reg181) : $unsigned(forvar260))}) | reg216[(3'h6):(3'h4)]);
              reg354 = (reg344 + ((8'hac) ^ $unsigned((!$signed((8'ha9))))));
              reg355 = $signed(({(reg275 != $unsigned(forvar346))} <= forvar254));
            end
          for (forvar356 = (1'h0); (forvar356 < (2'h2)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 = (~|wire174);
              reg358 <= $unsigned(reg181);
              reg359 = $signed(reg234[(3'h5):(3'h4)]);
              reg360 = $signed("N4a220");
              reg361 = ($unsigned((~&$signed((&(8'ha4))))) ?
                  forvar337[(3'h4):(2'h2)] : $unsigned(reg259[(4'hb):(3'h6)]));
            end
        end
      reg362 = ($unsigned($signed(forvar260[(1'h0):(1'h0)])) < ($signed(reg272[(2'h2):(1'h1)]) ?
          ($unsigned((8'hb5)) ?
              (((8'ha9) ? reg345 : reg216) <= (forvar319 ?
                  reg239 : reg211)) : (~^$unsigned(forvar351))) : $signed((~|(forvar309 ?
              reg181 : forvar207)))));
      reg363 <= reg354[(4'he):(2'h3)];
    end
  assign wire364 = $signed(reg261[(1'h0):(1'h0)]);
  assign wire365 = $unsigned(reg318[(2'h2):(1'h1)]);
  assign wire366 = (8'had);
  assign wire367 = {$signed({(forvar182 >= (-reg293)), (~^(+reg250))})};
  assign wire368 = (wire178 ^ ((&$unsigned({reg324})) ? (+reg323) : wire177));
  assign wire369 = ((^~{(reg253 ?
                           $unsigned(reg226) : ((8'ha6) ?
                               reg211 : reg212))}) != (|$unsigned($unsigned((reg320 ?
                       (8'hb4) : reg324)))));
  assign wire370 = forvar337[(2'h3):(2'h3)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module33
#( parameter param98 = (^(+(~(((8'ha0) ^ (8'hb8)) ? {(7'h41), (8'hb2)} : ((7'h42) ? (8'ha3) : (8'h9c)))))) )
(y, clk, wire37, wire36, wire35, wire34);
  output wire [(32'h2a0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire37;
  input wire [(4'hf):(1'h0)] wire36;
  input wire signed [(5'h11):(1'h0)] wire35;
  input wire [(3'h4):(1'h0)] wire34;
  reg signed [(4'h8):(1'h0)] reg97 = (1'h0);
  reg [(5'h14):(1'h0)] forvar96 = (1'h0);
  reg [(2'h2):(1'h0)] reg95 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar94 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg93 = (1'h0);
  reg [(3'h7):(1'h0)] reg92 = (1'h0);
  reg [(3'h7):(1'h0)] reg91 = (1'h0);
  reg [(4'he):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar87 = (1'h0);
  reg [(4'h8):(1'h0)] reg86 = (1'h0);
  reg [(4'h8):(1'h0)] reg85 = (1'h0);
  reg [(5'h11):(1'h0)] forvar84 = (1'h0);
  reg [(3'h5):(1'h0)] reg83 = (1'h0);
  reg [(4'ha):(1'h0)] reg82 = (1'h0);
  reg [(5'h15):(1'h0)] forvar81 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar80 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg79 = (1'h0);
  reg [(5'h10):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar77 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg76 = (1'h0);
  reg [(5'h12):(1'h0)] forvar75 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar73 = (1'h0);
  reg [(4'hf):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg71 = (1'h0);
  reg [(5'h13):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg68 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar67 = (1'h0);
  reg [(4'he):(1'h0)] reg66 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar64 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg61 = (1'h0);
  reg [(2'h3):(1'h0)] forvar60 = (1'h0);
  reg [(3'h5):(1'h0)] forvar59 = (1'h0);
  reg [(4'h8):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg57 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg56 = (1'h0);
  reg [(5'h13):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg54 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg53 = (1'h0);
  reg [(3'h5):(1'h0)] reg52 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar51 = (1'h0);
  reg [(3'h6):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg49 = (1'h0);
  reg [(4'ha):(1'h0)] reg48 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg47 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg46 = (1'h0);
  reg [(4'hb):(1'h0)] reg45 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg44 = (1'h0);
  reg [(3'h6):(1'h0)] forvar43 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar42 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire41;
  wire signed [(4'hd):(1'h0)] wire40;
  reg [(5'h14):(1'h0)] reg39 = (1'h0);
  reg signed [(4'he):(1'h0)] reg38 = (1'h0);
  assign y = {reg97,
                 forvar96,
                 reg95,
                 forvar94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 forvar87,
                 reg86,
                 reg85,
                 forvar84,
                 reg83,
                 reg82,
                 forvar81,
                 forvar80,
                 reg79,
                 reg78,
                 forvar77,
                 reg76,
                 forvar75,
                 reg74,
                 forvar73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 forvar67,
                 reg66,
                 reg65,
                 forvar64,
                 reg63,
                 reg62,
                 reg61,
                 forvar60,
                 forvar59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 forvar51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 forvar43,
                 forvar42,
                 wire41,
                 wire40,
                 reg39,
                 reg38,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg38 = wire37;
      reg39 <= wire34[(1'h1):(1'h1)];
    end
  assign wire40 = wire37[(3'h5):(1'h1)];
  assign wire41 = ((wire40 ?
                          ($unsigned(reg39) ?
                              $signed($signed(wire35)) : reg39[(3'h6):(3'h4)]) : reg38) ?
                      wire37 : (8'hb5));
  always
    @(posedge clk) begin
      for (forvar42 = (1'h0); (forvar42 < (1'h1)); forvar42 = (forvar42 + (1'h1)))
        begin
          for (forvar43 = (1'h0); (forvar43 < (1'h0)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg44 <= $unsigned($signed(wire37));
              reg45 = (8'hae);
              reg46 = $unsigned($signed($unsigned(((reg39 || reg44) ?
                  $signed(reg45) : reg39))));
            end
          reg47 = $unsigned((&($signed($unsigned(forvar43)) && ($signed(wire36) ?
              (-wire36) : (reg44 ? wire35 : reg38)))));
        end
    end
  always
    @(posedge clk) begin
      reg48 <= (~&$unsigned((((wire35 >> (8'ha4)) ?
              ((8'ha1) ? forvar42 : reg44) : forvar43) ?
          wire41 : wire41[(1'h1):(1'h1)])));
      reg49 <= wire40[(4'h9):(1'h0)];
      reg50 = ($unsigned((^~(+$signed(wire36)))) && ($unsigned({{(8'haf)},
          (wire34 ?
              wire37 : reg44)}) + (wire40[(1'h0):(1'h0)] >>> ($signed(forvar42) != reg45))));
      if ((wire36 ? (8'haa) : $unsigned(reg39[(1'h0):(1'h0)])))
        begin
          for (forvar51 = (1'h0); (forvar51 < (3'h4)); forvar51 = (forvar51 + (1'h1)))
            begin
              reg52 <= (wire36 ?
                  (($unsigned($signed(reg49)) >>> $unsigned((~|forvar42))) ?
                      $unsigned($signed(forvar51[(3'h6):(3'h4)])) : wire36[(3'h7):(2'h3)]) : (wire36 > $signed((~&forvar43))));
              reg53 <= reg49;
              reg54 = (8'hae);
              reg55 <= (($unsigned(((reg39 ?
                  wire36 : wire37) <<< reg45[(1'h1):(1'h1)])) + reg38[(4'hd):(4'ha)]) <= ({(!reg44)} ?
                  wire35 : $signed($signed(reg47))));
            end
        end
      else
        begin
          for (forvar51 = (1'h0); (forvar51 < (2'h2)); forvar51 = (forvar51 + (1'h1)))
            begin
              reg52 = ($unsigned($unsigned({(reg44 <= reg52)})) ^ reg49[(3'h5):(2'h3)]);
              reg53 = reg39[(3'h7):(1'h0)];
            end
          if (reg50[(3'h6):(1'h1)])
            begin
              reg54 <= reg46[(2'h2):(1'h0)];
              reg55 = (((^~(-reg45[(4'h9):(3'h5)])) ?
                      ($signed({(8'h9c)}) ?
                          reg53[(1'h1):(1'h0)] : (8'ha6)) : (~&(-(forvar43 ?
                          wire35 : wire40)))) ?
                  {(8'hb0),
                      $unsigned($unsigned(reg44[(3'h4):(2'h3)]))} : ((8'hb3) > reg50[(3'h5):(1'h0)]));
              reg56 <= reg54;
              reg57 <= (+(((&(reg47 > reg56)) != forvar51[(1'h0):(1'h0)]) >> reg47[(2'h2):(2'h2)]));
            end
          else
            begin
              reg54 <= $signed((({forvar42[(1'h1):(1'h1)]} ?
                      (wire37 ? $unsigned(reg54) : (+reg48)) : (reg44 * (reg48 ?
                          (8'hab) : (8'hba)))) ?
                  (^~((forvar42 ? forvar51 : forvar43) ?
                      (reg39 ^~ wire36) : (reg49 | wire35))) : wire34));
              reg55 = ((~&$unsigned($signed(((8'hb9) ?
                  reg44 : wire35)))) >= (wire35 ?
                  (((^reg45) * (reg50 && wire40)) ?
                      forvar43[(2'h3):(1'h0)] : ("BQ0Iv" - {reg47})) : (((reg46 ~^ (8'had)) ?
                      (reg44 ^~ reg48) : $signed((8'ha9))) > $unsigned({reg50,
                      forvar43}))));
              reg56 <= $unsigned((^~reg47[(1'h0):(1'h0)]));
              reg57 <= (reg48 ?
                  $unsigned((~^$unsigned((|reg52)))) : $signed(reg53[(1'h1):(1'h1)]));
            end
          reg58 = (^~$signed(($unsigned("GyRX") >>> (7'h41))));
        end
      for (forvar59 = (1'h0); (forvar59 < (2'h2)); forvar59 = (forvar59 + (1'h1)))
        begin
          for (forvar60 = (1'h0); (forvar60 < (1'h0)); forvar60 = (forvar60 + (1'h1)))
            begin
              reg61 <= $unsigned(forvar59[(1'h1):(1'h1)]);
              reg62 = (~|($unsigned(reg55) ^ (+(7'h44))));
              reg63 = ($unsigned(((~&"DbnHoGPJx") ?
                  $signed($signed((8'hbd))) : $unsigned(forvar59[(2'h2):(2'h2)]))) || {$unsigned("m")});
            end
          for (forvar64 = (1'h0); (forvar64 < (1'h1)); forvar64 = (forvar64 + (1'h1)))
            begin
              reg65 <= forvar60[(1'h0):(1'h0)];
              reg66 <= reg44;
            end
          for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= (({forvar42[(3'h7):(3'h5)],
                          $unsigned($unsigned(reg54))} ?
                      (reg52 <= ((reg38 ? (8'ha0) : (7'h43)) ?
                          {wire36,
                              (8'h9f)} : $signed(reg44))) : (-$signed((&(8'h9c))))) ?
                  (~^reg52[(1'h0):(1'h0)]) : $unsigned((8'hb6)));
              reg69 = (+$signed(wire36[(2'h2):(2'h2)]));
              reg70 = forvar43[(1'h1):(1'h0)];
              reg71 = reg61;
              reg72 = reg62[(3'h6):(3'h6)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar73 = (1'h0); (forvar73 < (3'h4)); forvar73 = (forvar73 + (1'h1)))
        begin
          reg74 <= (reg44[(4'h9):(3'h6)] << (+((~(|(8'hb8))) <<< wire36)));
        end
      for (forvar75 = (1'h0); (forvar75 < (3'h4)); forvar75 = (forvar75 + (1'h1)))
        begin
          reg76 <= reg62[(4'ha):(2'h2)];
          for (forvar77 = (1'h0); (forvar77 < (1'h1)); forvar77 = (forvar77 + (1'h1)))
            begin
              reg78 = $signed((^("ZJ1VYr8UhMMXyZ5" ?
                  reg50[(2'h3):(2'h2)] : wire36[(4'ha):(1'h1)])));
              reg79 = reg65;
            end
        end
      for (forvar80 = (1'h0); (forvar80 < (2'h2)); forvar80 = (forvar80 + (1'h1)))
        begin
          for (forvar81 = (1'h0); (forvar81 < (2'h3)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 <= ((~^reg44) ?
                  $unsigned("PeeUdd5VcaiT7W") : (!$unsigned(forvar64)));
              reg83 = ((reg76 ?
                  $signed((~&reg63)) : $signed((-(reg65 == reg71)))) + ($signed("LlkOg7Ww4XpREqm4uJpd") ?
                  ((^~reg56[(2'h2):(1'h1)]) <<< forvar77) : (^{reg62,
                      (forvar42 >= reg46)})));
            end
          for (forvar84 = (1'h0); (forvar84 < (1'h1)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 <= {{$unsigned((8'ha5))},
                  (($unsigned((wire41 ? reg52 : (8'ha4))) ?
                          (^reg48) : (8'hb4)) ?
                      ($signed((forvar59 >> (8'hb9))) ?
                          $signed($unsigned(forvar67)) : $unsigned({reg69})) : reg72[(3'h4):(1'h1)])};
            end
          reg86 <= {$unsigned({reg50, reg72[(1'h0):(1'h0)]})};
        end
      for (forvar87 = (1'h0); (forvar87 < (3'h4)); forvar87 = (forvar87 + (1'h1)))
        begin
          if (reg46[(1'h0):(1'h0)])
            begin
              reg88 = (-$unsigned($unsigned(((^forvar81) >>> $signed(reg82)))));
              reg89 <= ((^(~$signed($signed((7'h43))))) < reg54);
              reg90 = $signed({$signed(reg61[(4'h8):(3'h5)])});
              reg91 = ((reg86 - reg79[(2'h3):(2'h3)]) ?
                  (~($signed(reg62) | (8'had))) : (wire37[(3'h6):(2'h3)] - (-reg46[(2'h2):(2'h2)])));
            end
          else
            begin
              reg88 = $unsigned((reg71 ? forvar80 : $unsigned(wire35)));
              reg89 <= $unsigned(reg38[(4'h8):(1'h0)]);
            end
          reg92 <= reg50[(3'h4):(1'h0)];
          reg93 <= $unsigned($unsigned(($signed((wire36 ?
              forvar81 : reg70)) * reg69)));
        end
      for (forvar94 = (1'h0); (forvar94 < (1'h0)); forvar94 = (forvar94 + (1'h1)))
        begin
          reg95 <= (8'hb0);
          for (forvar96 = (1'h0); (forvar96 < (1'h1)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 = $unsigned(((8'hb0) ?
                  $signed(reg52[(3'h4):(3'h4)]) : (!reg86[(1'h0):(1'h0)])));
            end
        end
    end
endmodule
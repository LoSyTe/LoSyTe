(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param554 = (((^(((7'h41) ? (8'ha3) : (8'hb8)) >= ((8'h9c) >>> (8'hb1)))) - (((8'hb0) <= ((8'h9d) * (7'h42))) ? (((8'hb5) ? (8'ha2) : (8'hbd)) >> {(8'hb2), (8'h9c)}) : (|((8'h9d) ? (8'hba) : (8'ha5))))) || ((^~(((8'hbc) ? (8'ha7) : (7'h42)) ? {(8'hb5)} : ((8'ha8) * (8'hb8)))) <<< (^(8'h9c)))))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h425):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire0;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire [(4'hb):(1'h0)] wire3;
  wire [(2'h2):(1'h0)] wire553;
  wire [(4'h8):(1'h0)] wire552;
  wire [(3'h5):(1'h0)] wire535;
  wire signed [(4'hd):(1'h0)] wire468;
  wire signed [(5'h12):(1'h0)] wire466;
  wire signed [(4'hf):(1'h0)] wire465;
  wire signed [(5'h13):(1'h0)] wire464;
  wire signed [(4'hd):(1'h0)] wire457;
  wire [(5'h14):(1'h0)] wire459;
  wire signed [(5'h14):(1'h0)] wire460;
  wire signed [(5'h11):(1'h0)] wire461;
  wire [(5'h14):(1'h0)] wire462;
  wire signed [(4'ha):(1'h0)] wire470;
  reg signed [(2'h3):(1'h0)] reg548 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg549 = (1'h0);
  reg [(3'h7):(1'h0)] reg545 = (1'h0);
  reg [(4'ha):(1'h0)] reg544 = (1'h0);
  reg [(2'h3):(1'h0)] reg543 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg541 = (1'h0);
  reg [(2'h3):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg537 = (1'h0);
  reg [(5'h13):(1'h0)] reg533 = (1'h0);
  reg [(4'h9):(1'h0)] reg532 = (1'h0);
  reg [(4'he):(1'h0)] reg531 = (1'h0);
  reg [(2'h3):(1'h0)] reg525 = (1'h0);
  reg [(3'h6):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg523 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg520 = (1'h0);
  reg [(5'h12):(1'h0)] reg518 = (1'h0);
  reg [(2'h3):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg513 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg511 = (1'h0);
  reg [(4'hc):(1'h0)] reg510 = (1'h0);
  reg [(3'h7):(1'h0)] reg508 = (1'h0);
  reg [(4'ha):(1'h0)] reg505 = (1'h0);
  reg [(4'he):(1'h0)] reg504 = (1'h0);
  reg [(2'h3):(1'h0)] reg502 = (1'h0);
  reg [(3'h5):(1'h0)] reg500 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg499 = (1'h0);
  reg [(2'h3):(1'h0)] reg498 = (1'h0);
  reg [(4'hf):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg496 = (1'h0);
  reg [(5'h10):(1'h0)] reg493 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg491 = (1'h0);
  reg [(5'h13):(1'h0)] reg490 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg488 = (1'h0);
  reg [(5'h15):(1'h0)] reg486 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg485 = (1'h0);
  reg [(4'hb):(1'h0)] reg481 = (1'h0);
  reg [(5'h10):(1'h0)] reg479 = (1'h0);
  reg [(4'he):(1'h0)] reg472 = (1'h0);
  reg [(4'h8):(1'h0)] reg477 = (1'h0);
  reg [(4'hf):(1'h0)] reg476 = (1'h0);
  reg [(4'h8):(1'h0)] reg475 = (1'h0);
  reg [(5'h11):(1'h0)] reg474 = (1'h0);
  reg [(4'hd):(1'h0)] reg473 = (1'h0);
  reg [(4'ha):(1'h0)] reg550 = (1'h0);
  reg [(5'h10):(1'h0)] forvar548 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg547 = (1'h0);
  reg [(4'hb):(1'h0)] reg546 = (1'h0);
  reg [(3'h5):(1'h0)] forvar542 = (1'h0);
  reg [(5'h14):(1'h0)] forvar540 = (1'h0);
  reg [(4'he):(1'h0)] forvar538 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar536 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg534 = (1'h0);
  reg [(4'h9):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar529 = (1'h0);
  reg [(4'hd):(1'h0)] forvar528 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg526 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg522 = (1'h0);
  reg [(4'h9):(1'h0)] reg521 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg517 = (1'h0);
  reg [(4'hc):(1'h0)] reg516 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar515 = (1'h0);
  reg [(4'h8):(1'h0)] reg512 = (1'h0);
  reg [(5'h11):(1'h0)] reg509 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar507 = (1'h0);
  reg [(4'hb):(1'h0)] reg506 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar503 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg501 = (1'h0);
  reg [(4'h9):(1'h0)] forvar495 = (1'h0);
  reg [(2'h2):(1'h0)] forvar494 = (1'h0);
  reg [(3'h7):(1'h0)] forvar492 = (1'h0);
  reg [(4'he):(1'h0)] forvar489 = (1'h0);
  reg [(4'he):(1'h0)] reg487 = (1'h0);
  reg [(5'h15):(1'h0)] reg484 = (1'h0);
  reg [(2'h3):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg480 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg478 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar472 = (1'h0);
  assign y = {wire553,
                 wire552,
                 wire535,
                 wire468,
                 wire466,
                 wire465,
                 wire464,
                 wire457,
                 wire459,
                 wire460,
                 wire461,
                 wire462,
                 wire470,
                 reg548,
                 reg551,
                 reg549,
                 reg545,
                 reg544,
                 reg543,
                 reg541,
                 reg539,
                 reg537,
                 reg533,
                 reg532,
                 reg531,
                 reg525,
                 reg524,
                 reg523,
                 reg520,
                 reg518,
                 reg514,
                 reg513,
                 reg511,
                 reg510,
                 reg508,
                 reg505,
                 reg504,
                 reg502,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg493,
                 reg491,
                 reg490,
                 reg488,
                 reg486,
                 reg485,
                 reg481,
                 reg479,
                 reg472,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg550,
                 forvar548,
                 reg547,
                 reg546,
                 forvar542,
                 forvar540,
                 forvar538,
                 forvar536,
                 reg534,
                 reg530,
                 forvar529,
                 forvar528,
                 reg527,
                 reg526,
                 reg522,
                 reg521,
                 forvar519,
                 reg517,
                 reg516,
                 forvar515,
                 reg512,
                 reg509,
                 forvar507,
                 reg506,
                 forvar503,
                 reg501,
                 forvar495,
                 forvar494,
                 forvar492,
                 forvar489,
                 reg487,
                 reg484,
                 reg483,
                 forvar482,
                 reg480,
                 reg478,
                 forvar472,
                 (1'h0)};
  module4 #() modinst458 (wire457, clk, wire0, wire3, wire1, wire2, (8'ha6));
  assign wire459 = "6cbPFfThZD82yAqP3pu";
  assign wire460 = $signed($unsigned(wire0[(4'he):(4'he)]));
  assign wire461 = $unsigned($signed($signed(((wire0 ? wire460 : wire3) ?
                       $unsigned(wire1) : (wire2 && (8'hb8))))));
  module157 #() modinst463 (wire462, clk, wire2, wire461, wire459, wire1, wire460);
  assign wire464 = {((8'hab) ~^ $unsigned($unsigned({wire2}))),
                       $unsigned((wire462[(4'hc):(4'hc)] ?
                           "HV75WqtTH01tgNs3oKVB" : wire457[(3'h4):(2'h3)]))};
  assign wire465 = wire461;
  module325 #() modinst467 (.clk(clk), .y(wire466), .wire327(wire459), .wire328(wire462), .wire326(wire2), .wire329(wire457));
  module4 #() modinst469 (wire468, clk, wire2, wire457, wire466, wire461, wire459);
  module11 #() modinst471 (.wire13(wire466), .wire12(wire465), .wire16(wire460), .y(wire470), .clk(clk), .wire15(wire468), .wire14(wire3));
  always
    @(posedge clk) begin
      if (wire465)
        begin
          for (forvar472 = (1'h0); (forvar472 < (2'h3)); forvar472 = (forvar472 + (1'h1)))
            begin
              reg473 <= wire461;
              reg474 <= wire462;
              reg475 <= wire1;
              reg476 <= $unsigned($signed(((~(wire0 && wire2)) | "3DJZM2wc9piyiDTbT4U1")));
              reg477 <= reg474[(4'hb):(3'h4)];
            end
        end
      else
        begin
          reg472 <= $signed(wire470);
          if (forvar472[(1'h0):(1'h0)])
            begin
              reg478 = (~&forvar472[(2'h2):(1'h1)]);
              reg479 <= $signed(reg475);
              reg480 = $unsigned(wire461[(4'hf):(4'hc)]);
            end
          else
            begin
              reg473 <= $signed(wire464);
              reg478 = (~($signed(reg479) ?
                  $unsigned(($unsigned((8'haa)) ?
                      {reg479,
                          wire466} : reg480[(2'h3):(1'h1)])) : ((^~reg472[(1'h0):(1'h0)]) ?
                      ($unsigned(reg479) ?
                          wire3 : (&(8'ha5))) : {(reg476 | wire461)})));
              reg479 <= wire1;
            end
          reg481 <= $unsigned((($unsigned(wire1) ?
              wire459[(2'h2):(1'h0)] : (reg473[(4'hd):(4'hc)] ?
                  (~reg478) : {forvar472})) <= $signed((-(+reg480)))));
          for (forvar482 = (1'h0); (forvar482 < (2'h3)); forvar482 = (forvar482 + (1'h1)))
            begin
              reg483 = (!$unsigned((((!wire470) | wire462[(5'h13):(3'h5)]) ~^ $signed("gAVhh68lWpsX"))));
              reg484 = ((~^wire461) ?
                  $unsigned(wire2) : $signed({((reg478 > (8'ha6)) ?
                          $unsigned(wire459) : reg481)}));
              reg485 <= $unsigned(forvar472[(1'h0):(1'h0)]);
              reg486 <= $unsigned(((({wire464, wire2} > (reg483 ?
                      reg485 : reg483)) ^~ wire464[(4'hd):(4'hd)]) ?
                  $unsigned((~$unsigned(reg484))) : wire3[(1'h1):(1'h1)]));
              reg487 = wire462;
            end
        end
      reg488 <= ((reg486[(3'h5):(1'h1)] + reg484) > {reg475});
      for (forvar489 = (1'h0); (forvar489 < (3'h4)); forvar489 = (forvar489 + (1'h1)))
        begin
          reg490 <= (7'h41);
          reg491 <= reg487;
        end
      for (forvar492 = (1'h0); (forvar492 < (1'h1)); forvar492 = (forvar492 + (1'h1)))
        begin
          reg493 <= ((~|reg475) ? reg491[(1'h0):(1'h0)] : (|(7'h43)));
        end
      for (forvar494 = (1'h0); (forvar494 < (1'h0)); forvar494 = (forvar494 + (1'h1)))
        begin
          for (forvar495 = (1'h0); (forvar495 < (3'h4)); forvar495 = (forvar495 + (1'h1)))
            begin
              reg496 <= $unsigned((reg479 ?
                  {{forvar472[(1'h1):(1'h0)]}} : forvar494[(1'h1):(1'h0)]));
              reg497 <= $unsigned($signed(($signed($signed(reg491)) >= (wire464 ?
                  $unsigned(wire462) : {wire457, forvar489}))));
              reg498 <= $signed($signed((|forvar495[(1'h1):(1'h0)])));
            end
          if ((~((reg488[(4'he):(4'h8)] ?
                  $signed((reg480 ? wire457 : wire2)) : "s5X") ?
              $signed($unsigned((wire2 * wire3))) : (-($unsigned(reg480) >= {reg483,
                  wire462})))))
            begin
              reg499 <= $signed((~^(($signed((8'hb9)) == {reg497}) >= $unsigned(wire0))));
              reg500 <= (((((8'ha6) ?
                  $signed(forvar492) : {(8'hac),
                      wire464}) || $unsigned($signed(forvar482))) ^~ ((!(&(8'hb1))) != $unsigned((reg496 ?
                  reg479 : reg475)))) > "h");
              reg501 = $signed($unsigned(($unsigned($signed(wire464)) ?
                  (^reg472) : {{forvar482}})));
              reg502 <= {(("lLt5it1xn" ?
                          reg472 : ($unsigned(forvar489) ?
                              wire465 : ((7'h41) >>> wire3))) ?
                      (reg473 ?
                          ((reg490 ^ reg481) ?
                              (^~reg479) : $unsigned((8'ha2))) : ($signed(reg493) == "GLneZ3dr7rZpFVJXN")) : $unsigned($signed({forvar472}))),
                  reg501};
            end
          else
            begin
              reg499 <= ({reg488} > $signed($signed((-(reg500 & reg486)))));
              reg500 <= forvar482[(3'h7):(1'h0)];
              reg501 = reg484;
            end
          for (forvar503 = (1'h0); (forvar503 < (3'h4)); forvar503 = (forvar503 + (1'h1)))
            begin
              reg504 <= "nFqZ";
            end
          reg505 <= (&reg498);
        end
    end
  always
    @(posedge clk) begin
      reg506 = $unsigned({$signed(reg481), (~&wire460[(4'hf):(1'h1)])});
      for (forvar507 = (1'h0); (forvar507 < (2'h2)); forvar507 = (forvar507 + (1'h1)))
        begin
          if (((^~reg505[(3'h4):(1'h0)]) ? wire460 : reg474[(4'ha):(3'h7)]))
            begin
              reg508 <= $signed(reg499[(3'h4):(1'h0)]);
              reg509 = $signed($signed($unsigned($unsigned(reg486))));
              reg510 <= reg472;
              reg511 <= reg491[(3'h7):(3'h5)];
            end
          else
            begin
              reg509 = $signed(((^~{$signed(reg474),
                  (reg511 ? (7'h44) : reg493)}) ^~ $unsigned("")));
              reg512 = ($signed({((!forvar507) ?
                      $unsigned(reg472) : (wire457 != (8'had)))}) + ("c2CI5pqfYa4DliD" ?
                  wire470[(4'h9):(4'h8)] : {reg490}));
              reg513 <= (($signed(($unsigned(reg512) ?
                  (reg474 ^ (8'hb0)) : $unsigned(reg499))) >= ($unsigned((&reg474)) <= (+(reg485 ~^ wire3)))) & $unsigned(($signed(reg486) ?
                  forvar507 : (~|wire464))));
            end
          reg514 <= $signed($unsigned(reg505[(4'h9):(3'h7)]));
        end
      for (forvar515 = (1'h0); (forvar515 < (2'h3)); forvar515 = (forvar515 + (1'h1)))
        begin
          if ($unsigned((8'h9e)))
            begin
              reg516 = {$unsigned((~&((wire462 >= (7'h41)) ?
                      wire2 : (wire461 ? wire457 : wire465))))};
              reg517 = reg475;
            end
          else
            begin
              reg516 = ("639" == $signed(wire2));
              reg518 <= $signed((reg516[(2'h3):(1'h0)] != (($signed((8'hab)) ?
                      reg493 : (8'hb6)) ?
                  $unsigned((^~reg476)) : $signed($unsigned(reg511)))));
            end
          for (forvar519 = (1'h0); (forvar519 < (2'h3)); forvar519 = (forvar519 + (1'h1)))
            begin
              reg520 <= wire457;
            end
          reg521 = wire459[(5'h12):(4'hf)];
          if ({reg486[(4'ha):(1'h1)]})
            begin
              reg522 = $unsigned($unsigned((&forvar519)));
              reg523 <= (~&reg518[(3'h7):(2'h2)]);
              reg524 <= (^(reg505[(3'h6):(3'h5)] ?
                  (($unsigned(reg521) == (reg502 <<< (8'hb8))) < reg481) : (($unsigned(reg520) ?
                          {reg496, reg508} : (~&reg485)) ?
                      $signed((^reg514)) : $signed(reg504))));
              reg525 <= ($signed({(^~$unsigned(reg513)),
                      (&((7'h44) ? forvar507 : reg510))}) ?
                  ($unsigned(forvar515[(2'h2):(1'h1)]) ?
                      {((reg518 ^~ reg510) ?
                              {reg481, wire465} : reg472)} : (^$signed({(8'hac),
                          wire457}))) : "4MAuHGB1KD13bt3");
            end
          else
            begin
              reg522 = $signed((|((!$signed(wire1)) ?
                  wire457[(3'h4):(2'h3)] : $unsigned((^~reg510)))));
              reg526 = reg516[(4'hc):(4'hc)];
              reg527 = reg518;
            end
        end
      for (forvar528 = (1'h0); (forvar528 < (2'h2)); forvar528 = (forvar528 + (1'h1)))
        begin
          for (forvar529 = (1'h0); (forvar529 < (2'h3)); forvar529 = (forvar529 + (1'h1)))
            begin
              reg530 = ({wire1, reg514[(1'h0):(1'h0)]} ?
                  (((&"UcgHJRkekvXAcwTqaCq") * reg518[(4'h8):(3'h4)]) >>> (8'ha3)) : $signed((~wire3[(4'ha):(1'h0)])));
              reg531 <= reg504[(1'h1):(1'h0)];
              reg532 <= (~&reg510);
              reg533 <= reg512;
            end
        end
      reg534 = reg512[(4'h8):(1'h0)];
    end
  assign wire535 = (~|$signed(reg474));
  always
    @(posedge clk) begin
      for (forvar536 = (1'h0); (forvar536 < (2'h3)); forvar536 = (forvar536 + (1'h1)))
        begin
          reg537 <= reg502;
        end
      for (forvar538 = (1'h0); (forvar538 < (2'h2)); forvar538 = (forvar538 + (1'h1)))
        begin
          reg539 <= (~&$signed({(((8'ha0) && reg505) - (reg514 ?
                  wire535 : reg497)),
              reg477[(1'h1):(1'h0)]}));
        end
      for (forvar540 = (1'h0); (forvar540 < (1'h1)); forvar540 = (forvar540 + (1'h1)))
        begin
          reg541 <= (^reg476[(4'hf):(4'ha)]);
          for (forvar542 = (1'h0); (forvar542 < (1'h0)); forvar542 = (forvar542 + (1'h1)))
            begin
              reg543 <= (!(~($unsigned((reg532 ?
                  wire459 : reg500)) > reg493[(4'h8):(3'h5)])));
              reg544 <= $signed((((wire462[(5'h13):(1'h1)] ?
                  $unsigned(reg541) : $unsigned(reg525)) >>> $unsigned((reg539 ^~ wire0))) >= (&(8'h9f))));
              reg545 <= (~|(^$signed(reg524[(2'h3):(2'h3)])));
              reg546 = $unsigned(forvar540);
              reg547 = {({$unsigned((^~reg533)),
                      reg472} || ((^~$unsigned(wire457)) ?
                      reg520 : (~&(8'hb4))))};
            end
        end
      if ((8'had))
        begin
          for (forvar548 = (1'h0); (forvar548 < (2'h3)); forvar548 = (forvar548 + (1'h1)))
            begin
              reg549 <= reg524[(3'h4):(1'h0)];
              reg550 = ((~|$signed(({reg549, wire535} <= $signed(reg485)))) ?
                  $unsigned(wire466[(3'h4):(3'h4)]) : $signed(wire468[(4'h8):(3'h5)]));
            end
          reg551 <= (forvar540 * (wire466 ^~ reg511[(1'h1):(1'h1)]));
        end
      else
        begin
          reg548 <= reg537;
          reg549 <= reg475;
        end
    end
  assign wire552 = $unsigned((&{$unsigned((reg473 || reg539)),
                       {$unsigned((7'h41))}}));
  assign wire553 = reg518;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4  (y, clk, wire5, wire6, wire7, wire8, wire9);
  output wire [(32'h640):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire5;
  input wire [(3'h6):(1'h0)] wire6;
  input wire [(5'h11):(1'h0)] wire7;
  input wire signed [(5'h11):(1'h0)] wire8;
  input wire signed [(5'h14):(1'h0)] wire9;
  wire [(4'h9):(1'h0)] wire386;
  wire signed [(5'h14):(1'h0)] wire371;
  wire signed [(5'h12):(1'h0)] wire341;
  wire signed [(4'hc):(1'h0)] wire324;
  wire signed [(4'he):(1'h0)] wire323;
  wire [(4'hd):(1'h0)] wire322;
  wire [(4'hf):(1'h0)] wire321;
  wire [(5'h15):(1'h0)] wire320;
  wire [(4'hc):(1'h0)] wire151;
  wire [(5'h11):(1'h0)] wire133;
  wire signed [(5'h13):(1'h0)] wire10;
  wire signed [(4'hd):(1'h0)] wire131;
  wire signed [(5'h11):(1'h0)] wire153;
  wire [(4'hf):(1'h0)] wire154;
  wire signed [(4'hf):(1'h0)] wire155;
  wire [(4'h8):(1'h0)] wire156;
  wire signed [(5'h10):(1'h0)] wire318;
  reg [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(5'h11):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg451 = (1'h0);
  reg [(2'h2):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg446 = (1'h0);
  reg [(5'h10):(1'h0)] reg444 = (1'h0);
  reg [(3'h5):(1'h0)] reg440 = (1'h0);
  reg signed [(4'he):(1'h0)] reg439 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg438 = (1'h0);
  reg [(4'hb):(1'h0)] reg436 = (1'h0);
  reg [(4'hb):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg431 = (1'h0);
  reg [(4'hd):(1'h0)] reg430 = (1'h0);
  reg [(3'h5):(1'h0)] reg427 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg422 = (1'h0);
  reg [(4'hd):(1'h0)] reg419 = (1'h0);
  reg [(3'h6):(1'h0)] reg415 = (1'h0);
  reg [(2'h3):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg414 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg409 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg407 = (1'h0);
  reg [(5'h11):(1'h0)] reg406 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg404 = (1'h0);
  reg [(3'h4):(1'h0)] reg402 = (1'h0);
  reg [(5'h14):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg398 = (1'h0);
  reg [(2'h3):(1'h0)] reg397 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg395 = (1'h0);
  reg [(4'hf):(1'h0)] reg393 = (1'h0);
  reg [(3'h6):(1'h0)] reg392 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg391 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg389 = (1'h0);
  reg [(2'h3):(1'h0)] reg388 = (1'h0);
  reg [(4'ha):(1'h0)] reg383 = (1'h0);
  reg [(3'h4):(1'h0)] reg380 = (1'h0);
  reg [(4'ha):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] reg373 = (1'h0);
  reg [(4'ha):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg [(5'h11):(1'h0)] reg368 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg367 = (1'h0);
  reg [(4'he):(1'h0)] reg366 = (1'h0);
  reg [(4'hb):(1'h0)] reg365 = (1'h0);
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg361 = (1'h0);
  reg signed [(4'he):(1'h0)] reg360 = (1'h0);
  reg [(5'h10):(1'h0)] reg359 = (1'h0);
  reg [(4'h9):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg350 = (1'h0);
  reg [(4'hb):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg352 = (1'h0);
  reg [(5'h12):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg343 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg454 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg450 = (1'h0);
  reg [(3'h5):(1'h0)] forvar449 = (1'h0);
  reg [(5'h12):(1'h0)] reg447 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar441 = (1'h0);
  reg [(2'h2):(1'h0)] reg445 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg442 = (1'h0);
  reg [(4'ha):(1'h0)] reg441 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg437 = (1'h0);
  reg [(2'h3):(1'h0)] reg435 = (1'h0);
  reg [(4'ha):(1'h0)] forvar433 = (1'h0);
  reg [(4'hb):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg429 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar428 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg423 = (1'h0);
  reg [(3'h4):(1'h0)] forvar421 = (1'h0);
  reg [(3'h7):(1'h0)] reg420 = (1'h0);
  reg [(4'hd):(1'h0)] forvar418 = (1'h0);
  reg [(3'h6):(1'h0)] forvar414 = (1'h0);
  reg [(4'hc):(1'h0)] reg417 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar415 = (1'h0);
  reg [(4'h8):(1'h0)] reg413 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg405 = (1'h0);
  reg signed [(4'he):(1'h0)] reg403 = (1'h0);
  reg [(5'h11):(1'h0)] reg400 = (1'h0);
  reg [(3'h4):(1'h0)] forvar393 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg396 = (1'h0);
  reg [(4'ha):(1'h0)] reg394 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg390 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar387 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg385 = (1'h0);
  reg [(5'h14):(1'h0)] reg384 = (1'h0);
  reg [(4'he):(1'h0)] reg382 = (1'h0);
  reg [(4'he):(1'h0)] forvar381 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg379 = (1'h0);
  reg [(4'ha):(1'h0)] reg377 = (1'h0);
  reg [(4'hc):(1'h0)] reg376 = (1'h0);
  reg [(4'hd):(1'h0)] reg375 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar374 = (1'h0);
  reg [(4'hf):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg369 = (1'h0);
  reg [(2'h2):(1'h0)] forvar363 = (1'h0);
  reg [(4'ha):(1'h0)] reg362 = (1'h0);
  reg [(5'h13):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar357 = (1'h0);
  reg [(5'h14):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg353 = (1'h0);
  reg [(4'hb):(1'h0)] forvar350 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar346 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg345 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg344 = (1'h0);
  assign y = {wire386,
                 wire371,
                 wire341,
                 wire324,
                 wire323,
                 wire322,
                 wire321,
                 wire320,
                 wire151,
                 wire133,
                 wire10,
                 wire131,
                 wire153,
                 wire154,
                 wire155,
                 wire156,
                 wire318,
                 reg456,
                 reg455,
                 reg452,
                 reg451,
                 reg448,
                 reg446,
                 reg444,
                 reg440,
                 reg439,
                 reg438,
                 reg436,
                 reg434,
                 reg431,
                 reg430,
                 reg427,
                 reg426,
                 reg425,
                 reg422,
                 reg419,
                 reg415,
                 reg416,
                 reg414,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg404,
                 reg402,
                 reg401,
                 reg399,
                 reg398,
                 reg397,
                 reg395,
                 reg393,
                 reg392,
                 reg391,
                 reg389,
                 reg388,
                 reg383,
                 reg380,
                 reg378,
                 reg373,
                 reg372,
                 reg370,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg361,
                 reg360,
                 reg359,
                 reg356,
                 reg350,
                 reg355,
                 reg352,
                 reg351,
                 reg347,
                 reg343,
                 reg454,
                 reg453,
                 reg450,
                 forvar449,
                 reg447,
                 forvar441,
                 reg445,
                 reg443,
                 reg442,
                 reg441,
                 reg437,
                 reg435,
                 forvar433,
                 reg432,
                 reg429,
                 forvar428,
                 reg424,
                 reg423,
                 forvar421,
                 reg420,
                 forvar418,
                 forvar414,
                 reg417,
                 forvar415,
                 reg413,
                 reg412,
                 reg411,
                 reg405,
                 reg403,
                 reg400,
                 forvar393,
                 reg396,
                 reg394,
                 reg390,
                 forvar387,
                 reg385,
                 reg384,
                 reg382,
                 forvar381,
                 reg379,
                 reg377,
                 reg376,
                 reg375,
                 forvar374,
                 reg357,
                 reg369,
                 forvar363,
                 reg362,
                 reg358,
                 forvar357,
                 reg354,
                 reg353,
                 forvar350,
                 reg349,
                 reg348,
                 forvar346,
                 reg345,
                 reg344,
                 (1'h0)};
  assign wire10 = "Q9F8kPe4iuN3";
  module11 #() modinst132 (.y(wire131), .wire16(wire9), .wire14(wire5), .wire12(wire7), .wire13(wire10), .clk(clk), .wire15(wire8));
  assign wire133 = ((+(^~((wire8 ? wire9 : wire7) ?
                           {wire131} : (wire9 ? wire10 : wire10)))) ?
                       ($unsigned(($unsigned(wire8) ?
                               "qgTcSub2ceSXO69hii8n" : $unsigned(wire9))) ?
                           (7'h44) : (~&$signed((wire7 || wire9)))) : wire5);
  module134 #() modinst152 (.wire138(wire9), .y(wire151), .wire135(wire10), .wire139(wire8), .wire137(wire133), .wire136(wire7), .clk(clk));
  assign wire153 = wire7[(5'h10):(1'h0)];
  assign wire154 = $signed("FPl7Lxl8puxQ2Bf");
  assign wire155 = (wire131[(2'h3):(1'h1)] ?
                       $unsigned($unsigned((~&wire7[(1'h1):(1'h0)]))) : (|(~|({wire7} ?
                           wire9 : (-(8'hb6))))));
  assign wire156 = {wire10, (^(wire154[(4'h8):(3'h4)] >> wire151))};
  module157 #() modinst319 (.y(wire318), .wire158(wire153), .clk(clk), .wire161(wire155), .wire159(wire133), .wire162(wire9), .wire160(wire151));
  assign wire320 = (wire6 ?
                       (wire156[(3'h7):(1'h0)] ?
                           (-($unsigned(wire8) ?
                               $unsigned((8'hb1)) : $signed((8'hac)))) : wire9) : wire155[(4'hc):(1'h1)]);
  assign wire321 = $signed((^~(+{wire133[(3'h5):(3'h4)]})));
  assign wire322 = $signed($unsigned(($unsigned($unsigned(wire9)) ?
                       {(~&(8'ha0)),
                           ((8'hb5) ? wire318 : wire10)} : ($signed(wire320) ?
                           $unsigned(wire156) : $signed(wire321)))));
  assign wire323 = (wire7[(4'ha):(4'ha)] ?
                       (!(wire156[(3'h5):(1'h1)] * wire133)) : ($unsigned(wire320[(3'h7):(2'h2)]) * (&$unsigned({wire10,
                           wire5}))));
  assign wire324 = {$signed((~^({wire9} ^~ (^~wire155))))};
  module325 #() modinst342 (wire341, clk, wire324, wire7, wire155, wire5);
  always
    @(posedge clk) begin
      reg343 <= ((wire7[(3'h7):(2'h2)] ?
          (~(~&wire9)) : {(^~wire8[(5'h10):(1'h0)])}) >> wire154[(4'hb):(3'h6)]);
      reg344 = (^~(^~$signed(((wire6 ? wire9 : wire323) >= (~wire155)))));
      reg345 = ((8'hbe) ?
          (($signed(reg344[(4'h9):(3'h5)]) | (-$unsigned(wire320))) >>> wire151) : (&($signed({wire322,
                  wire10}) ?
              $unsigned((-wire153)) : (7'h44))));
      if ((~(($signed(wire322[(3'h6):(1'h1)]) ? "QgW" : $signed((~&reg343))) ?
          (reg343 ? wire154[(4'h9):(2'h2)] : $unsigned(wire341)) : {wire151})))
        begin
          for (forvar346 = (1'h0); (forvar346 < (1'h0)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 <= (~^($signed($unsigned(wire131)) <<< $unsigned(wire322[(4'hc):(2'h3)])));
              reg348 = wire156;
            end
          reg349 = wire324;
          for (forvar350 = (1'h0); (forvar350 < (3'h4)); forvar350 = (forvar350 + (1'h1)))
            begin
              reg351 <= wire318;
              reg352 <= (wire5[(5'h12):(2'h2)] >>> $signed(reg351));
              reg353 = wire318[(4'h8):(3'h7)];
              reg354 = ($unsigned(wire156) == wire154);
              reg355 <= (&($signed(((reg345 <<< wire8) ?
                      $signed(reg345) : $unsigned(wire318))) ?
                  (wire5[(4'hb):(2'h3)] * $signed((forvar350 ?
                      reg353 : forvar346))) : {{(wire321 != wire133),
                          $signed(wire155)},
                      wire7[(4'he):(4'h9)]}));
            end
        end
      else
        begin
          for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 <= ($signed(wire323[(4'hc):(4'h9)]) << (!reg355));
              reg348 = ("8p" && reg351);
              reg350 <= {$signed((|({wire133, (8'hbf)} || (wire324 ?
                      reg351 : wire320)))),
                  $unsigned((~(~|(forvar346 ? reg352 : forvar350))))};
              reg351 <= ("UysbECZZ3" ?
                  $unsigned(wire6) : (reg352 ?
                      (|(~$signed(wire321))) : (^~((wire153 ?
                              reg345 : (7'h44)) ?
                          $unsigned(wire153) : (wire156 > (8'hb3))))));
              reg352 <= $signed($unsigned($signed(("8BpuN7A" || $unsigned(wire5)))));
            end
          reg355 <= $unsigned($unsigned({(wire341[(4'h9):(3'h7)] ?
                  $unsigned(wire10) : wire131)}));
        end
    end
  always
    @(posedge clk) begin
      if (wire10)
        begin
          reg356 <= reg352[(5'h11):(3'h5)];
          for (forvar357 = (1'h0); (forvar357 < (1'h1)); forvar357 = (forvar357 + (1'h1)))
            begin
              reg358 = (wire320[(3'h7):(3'h7)] < ($unsigned($unsigned($signed(reg351))) ?
                  ((~(reg343 < reg356)) ?
                      {wire7,
                          ((8'hb4) ~^ forvar357)} : $signed($unsigned(reg343))) : (^~$unsigned($unsigned(wire7)))));
              reg359 <= wire6;
              reg360 <= (wire154 - "mhu");
              reg361 <= wire318[(1'h0):(1'h0)];
            end
          reg362 = $unsigned((wire8 > $signed(((reg343 ?
              (7'h42) : wire7) && $unsigned(wire131)))));
          for (forvar363 = (1'h0); (forvar363 < (2'h2)); forvar363 = (forvar363 + (1'h1)))
            begin
              reg364 <= ({$signed($signed({reg352, wire133})),
                      (($signed(wire155) ? (~|wire8) : (|(8'hab))) >> wire9)} ?
                  ($unsigned(((wire322 ? reg362 : wire322) < wire133)) ?
                      $signed($unsigned((~|reg350))) : ($unsigned((wire321 <= reg352)) || $signed({wire154}))) : (^~reg361));
              reg365 <= "GLUZw9H";
              reg366 <= ((((reg359[(2'h2):(1'h1)] ?
                      wire154[(2'h3):(2'h3)] : (~|wire324)) <<< {wire7,
                      reg364[(3'h5):(3'h5)]}) ?
                  (8'hb9) : (-$signed((~^reg361)))) || ((7'h42) < (&wire8)));
              reg367 <= wire341[(2'h2):(1'h1)];
              reg368 <= reg360;
            end
          reg369 = wire6[(1'h1):(1'h0)];
        end
      else
        begin
          reg357 = $unsigned(reg361);
          reg358 = reg355;
          reg362 = wire10[(5'h12):(4'hd)];
        end
      reg370 <= $unsigned((reg369 + ($signed((reg343 ?
          reg360 : reg365)) - wire320)));
    end
  assign wire371 = (-$signed($unsigned($unsigned(reg360[(4'h8):(3'h4)]))));
  always
    @(posedge clk) begin
      reg372 <= ((~|$unsigned($unsigned($unsigned(reg355)))) ?
          (wire153[(2'h3):(1'h1)] || $unsigned(reg359[(3'h5):(1'h0)])) : $signed((($signed(wire318) <= (~wire153)) != {wire10})));
      reg373 <= (+reg350);
      for (forvar374 = (1'h0); (forvar374 < (2'h2)); forvar374 = (forvar374 + (1'h1)))
        begin
          reg375 = (^~(8'hb4));
          if ({$unsigned(reg375[(3'h5):(3'h4)])})
            begin
              reg376 = (wire321[(4'h9):(1'h1)] ^ (~&(reg367[(3'h6):(3'h5)] ?
                  ((wire151 ?
                      reg366 : reg356) * wire131[(4'h8):(3'h4)]) : $unsigned(wire131[(1'h1):(1'h0)]))));
              reg377 = {((({wire318,
                      wire156} != wire6[(1'h0):(1'h0)]) != (8'ha7)) <= (!($unsigned(reg352) ?
                      wire8[(3'h6):(1'h1)] : $unsigned((8'hac))))),
                  $unsigned($unsigned("JO2AY1Ko"))};
            end
          else
            begin
              reg378 <= $signed($unsigned(reg366));
              reg379 = $unsigned($unsigned(({(~^reg351), (reg359 && (8'ha4))} ?
                  ((wire155 > reg377) ?
                      reg355 : (|reg355)) : (reg372[(4'h8):(3'h6)] ?
                      (wire156 || (8'h9f)) : reg347))));
            end
          reg380 <= $unsigned($unsigned(wire153));
        end
      for (forvar381 = (1'h0); (forvar381 < (1'h1)); forvar381 = (forvar381 + (1'h1)))
        begin
          if (wire324[(1'h0):(1'h0)])
            begin
              reg382 = {($unsigned(wire8[(4'hd):(1'h0)]) ?
                      (&reg350) : "buWrdod60QBZgO8RIxcX"),
                  {(-wire324[(3'h7):(3'h4)])}};
              reg383 <= {wire8};
              reg384 = $unsigned(wire155);
            end
          else
            begin
              reg382 = $unsigned((-$signed($unsigned({wire10, wire7}))));
              reg383 <= $signed($signed({(-((8'h9d) >= reg377))}));
              reg384 = reg375;
              reg385 = $signed(reg364);
            end
        end
    end
  assign wire386 = $signed(wire324);
  always
    @(posedge clk) begin
      for (forvar387 = (1'h0); (forvar387 < (2'h3)); forvar387 = (forvar387 + (1'h1)))
        begin
          if (wire8[(1'h1):(1'h0)])
            begin
              reg388 <= wire9[(2'h3):(2'h2)];
              reg389 <= reg378[(2'h2):(1'h1)];
              reg390 = wire8;
              reg391 <= reg359;
            end
          else
            begin
              reg388 <= ((reg351 > $signed(wire131[(4'hc):(3'h6)])) ?
                  ((!({(8'hae)} * $unsigned(reg366))) && {(~$signed((8'hb3))),
                      reg378}) : $signed($signed(reg350[(2'h2):(1'h0)])));
              reg389 <= {wire322[(4'hb):(4'ha)]};
            end
        end
      reg392 <= (8'ha3);
      if ((reg378 ^ (~&reg383)))
        begin
          if ({$unsigned(reg391),
              {(reg355[(2'h2):(2'h2)] ?
                      (wire7[(4'he):(4'ha)] ?
                          (wire154 & wire154) : $unsigned(forvar387)) : (+wire154)),
                  reg370[(4'h8):(4'h8)]}})
            begin
              reg393 <= (((&$signed(reg347)) * $signed($signed($signed(wire133)))) ^~ $unsigned(($unsigned((reg343 * reg351)) && (+((8'haf) - wire371)))));
              reg394 = (wire155 + ($signed({wire386[(4'h9):(4'h8)]}) + ("YY" ?
                  wire8[(1'h1):(1'h1)] : {(^~wire131)})));
            end
          else
            begin
              reg393 <= wire8[(1'h0):(1'h0)];
              reg395 <= (~|{"yuV6pz5wf"});
            end
          reg396 = $signed((|wire386[(3'h5):(3'h5)]));
        end
      else
        begin
          for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg395 <= ($unsigned($unsigned((8'haa))) ?
                  $signed(reg366) : $unsigned(({(reg360 == wire9), (8'hb5)} ?
                      $unsigned((^~reg343)) : (+$unsigned(reg388)))));
              reg397 <= (!(~wire131));
              reg398 <= (reg395 ? wire151 : (~|(8'h9e)));
            end
          if ($signed(reg380))
            begin
              reg399 <= ({$signed("uZ8LdhqJ9b"), $signed({(!reg366), reg392})} ?
                  wire386[(3'h4):(1'h0)] : $signed(reg347[(2'h2):(2'h2)]));
            end
          else
            begin
              reg400 = reg368[(3'h4):(1'h0)];
              reg401 <= (reg393[(4'hf):(4'hc)] ?
                  $unsigned(reg350[(4'hd):(2'h3)]) : $unsigned(wire318));
              reg402 <= $unsigned(($unsigned((&((8'hbd) << reg373))) ^ wire5[(4'hb):(4'h8)]));
              reg403 = (($signed(reg360[(4'h9):(3'h4)]) <= $unsigned(reg343[(4'hb):(3'h6)])) ?
                  $signed((wire154 >>> ($unsigned(wire8) ?
                      $signed(forvar387) : ((7'h41) ~^ reg391)))) : wire154);
              reg404 <= reg396;
            end
          if (forvar393[(3'h4):(2'h2)])
            begin
              reg405 = $unsigned($signed((^((reg390 == reg400) + (|wire386)))));
            end
          else
            begin
              reg406 <= $unsigned(wire318[(3'h5):(2'h3)]);
              reg407 <= $unsigned(({$unsigned(reg343[(2'h3):(2'h3)])} ?
                  (8'hbb) : (~|$signed((reg355 ? wire151 : reg356)))));
            end
          reg408 <= $unsigned($signed((8'had)));
          reg409 <= $signed(reg401);
        end
      if (wire156)
        begin
          reg410 <= (8'hb0);
          if (reg407)
            begin
              reg411 = $signed((!$signed((~|wire7))));
              reg412 = {{reg400[(1'h1):(1'h0)]}, reg410};
              reg413 = ((forvar387 || reg350[(4'hf):(3'h4)]) == reg400);
            end
          else
            begin
              reg414 <= ($signed(wire154) << (~^($signed(reg356) & reg413[(1'h0):(1'h0)])));
            end
          for (forvar415 = (1'h0); (forvar415 < (2'h3)); forvar415 = (forvar415 + (1'h1)))
            begin
              reg416 <= {({(wire10[(3'h6):(1'h0)] ?
                          wire371 : reg414)} <<< (~&(reg406 ?
                      reg378[(3'h5):(3'h4)] : (-wire386)))),
                  {(+($unsigned(reg359) != reg405)), wire321}};
            end
          reg417 = (((^~{(wire10 & reg395),
              $unsigned(reg396)}) != $signed($unsigned(reg373))) | ($signed(reg350) >>> reg389));
        end
      else
        begin
          if (($signed(reg416[(1'h1):(1'h0)]) ^ reg350))
            begin
              reg411 = $unsigned(($signed(reg409[(4'hb):(1'h0)]) ?
                  (~|(wire7[(4'hd):(4'h8)] ?
                      (!reg343) : (wire9 == reg352))) : (~^(wire10 > (~|wire322)))));
              reg412 = (+$unsigned($unsigned(reg398)));
              reg413 = wire7;
            end
          else
            begin
              reg410 <= (reg364 ?
                  $signed(wire320[(4'hf):(3'h7)]) : {$signed((reg392[(2'h3):(2'h3)] || "")),
                      $signed(reg403[(4'h9):(1'h1)])});
              reg411 = $unsigned(($signed(((wire386 | reg410) ?
                      (reg398 ? reg373 : wire341) : $unsigned((8'had)))) ?
                  reg360 : (($signed(reg360) - (^~reg394)) >= {(reg401 ?
                          reg372 : reg370),
                      (~|reg397)})));
            end
          for (forvar414 = (1'h0); (forvar414 < (2'h3)); forvar414 = (forvar414 + (1'h1)))
            begin
              reg415 <= ($unsigned(reg380[(1'h1):(1'h0)]) < (wire9 > reg416));
              reg417 = wire156[(4'h8):(2'h2)];
            end
        end
      for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
        begin
          reg419 <= $signed(reg364);
          reg420 = $unsigned($unsigned(((wire371[(4'h9):(3'h6)] * (~&reg373)) ?
              ((+forvar415) ^~ (reg356 ?
                  (8'had) : wire371)) : reg365[(1'h1):(1'h0)])));
          for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= "3kPZhSFsyIEh";
              reg423 = reg394;
              reg424 = reg366[(4'hd):(4'hb)];
              reg425 <= ($unsigned((reg350 ?
                  wire321[(4'ha):(4'h9)] : $unsigned($unsigned(reg372)))) + ((~|(!wire321)) <= (7'h44)));
              reg426 <= reg350[(4'he):(4'h9)];
            end
          reg427 <= $signed($unsigned(($signed(reg398[(4'hb):(4'h9)]) & (~&$unsigned(wire153)))));
          for (forvar428 = (1'h0); (forvar428 < (3'h4)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 = {reg351};
              reg430 <= ((~^(~{"hLC2"})) ?
                  $signed($signed($unsigned((reg392 ~^ reg400)))) : {$unsigned(reg391[(3'h6):(2'h2)]),
                      reg413});
              reg431 <= {wire156};
            end
        end
    end
  always
    @(posedge clk) begin
      reg432 = (reg361[(4'hc):(3'h6)] ?
          reg409[(4'hd):(2'h3)] : ({((~wire386) ?
                      $signed(reg343) : {reg359, reg370}),
                  reg370} ?
              reg364[(3'h7):(1'h0)] : wire154));
      if (($unsigned((~^{$signed(reg395)})) ?
          {(wire318[(2'h2):(1'h1)] ? (8'hab) : reg409[(3'h4):(2'h3)])} : wire5))
        begin
          for (forvar433 = (1'h0); (forvar433 < (2'h2)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= reg388;
              reg435 = (-reg368);
              reg436 <= reg380[(2'h2):(2'h2)];
              reg437 = $unsigned((reg391 & reg422[(3'h5):(3'h4)]));
            end
          reg438 <= (~|wire133[(3'h7):(3'h7)]);
          if ("0cu9k6nl7xsQ6x")
            begin
              reg439 <= (~(~&$unsigned(reg410)));
              reg440 <= (8'haa);
              reg441 = wire10;
            end
          else
            begin
              reg441 = wire318;
              reg442 = $signed((^(reg350 >= (8'ha9))));
              reg443 = wire154[(4'h8):(3'h7)];
              reg444 <= ($signed((^reg364)) >>> $signed($unsigned(((+reg367) ?
                  (reg425 << wire321) : (reg399 ^ (8'ha6))))));
            end
          reg445 = ((reg392[(2'h3):(2'h3)] >> (-reg416[(2'h2):(1'h1)])) ?
              ($unsigned($unsigned(wire151)) <<< ($unsigned({reg438, wire5}) ?
                  reg352 : reg392[(1'h0):(1'h0)])) : ($unsigned({wire7,
                      reg402}) ?
                  reg347[(3'h4):(3'h4)] : ($unsigned(reg364) ?
                      reg343 : $signed($signed(reg441)))));
          reg446 <= (&$unsigned(reg398[(4'hd):(3'h7)]));
        end
      else
        begin
          for (forvar433 = (1'h0); (forvar433 < (1'h0)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= $unsigned($signed($signed(reg366[(4'hc):(3'h7)])));
              reg436 <= {wire155[(3'h4):(2'h3)],
                  ($signed((~&{reg367})) ^~ $unsigned(((reg446 >>> (8'ha2)) ^~ (!reg445))))};
              reg438 <= $signed(reg439);
              reg439 <= ((!$signed(wire341[(4'h8):(3'h6)])) * $unsigned(reg380[(1'h1):(1'h1)]));
            end
          reg440 <= reg406;
          for (forvar441 = (1'h0); (forvar441 < (3'h4)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 = (&(!{reg437[(3'h6):(1'h1)], "Rwbk"}));
              reg444 <= wire7[(3'h6):(3'h4)];
              reg445 = (~wire9[(2'h2):(1'h0)]);
            end
          if ({$signed({$unsigned($signed(wire9))})})
            begin
              reg447 = ((~&($unsigned((reg415 && reg437)) ^ wire324)) || $signed(({(!reg437)} ?
                  (8'hac) : $unsigned($unsigned(wire322)))));
              reg448 <= reg350;
            end
          else
            begin
              reg447 = ((-$signed((-$signed(wire324)))) && (^($signed($signed((8'h9c))) ?
                  $unsigned((wire318 || (8'had))) : $unsigned($unsigned(wire5)))));
            end
        end
      if (wire318)
        begin
          for (forvar449 = (1'h0); (forvar449 < (2'h2)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 = reg445[(2'h2):(2'h2)];
              reg451 <= $unsigned((reg447[(2'h3):(2'h2)] ?
                  $unsigned((reg406 && wire322[(3'h5):(3'h4)])) : ((8'hb5) ~^ $unsigned({wire154,
                      reg425}))));
              reg452 <= ($signed($signed($signed({reg448,
                  (8'ha9)}))) < {reg450[(3'h4):(1'h1)]});
            end
        end
      else
        begin
          for (forvar449 = (1'h0); (forvar449 < (1'h0)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg451 <= (reg438 ?
                  (~((~|reg359[(2'h2):(1'h0)]) ?
                      {(reg351 ? reg356 : wire155),
                          (reg437 ?
                              (8'ha7) : wire9)} : $signed(reg446))) : $unsigned($signed($signed((8'ha7)))));
              reg452 <= $unsigned(((|wire320) < reg361));
              reg453 = $signed({(((&reg426) ? reg439 : $unsigned(reg422)) ?
                      reg370 : (wire324 ? wire371 : wire341)),
                  $signed($unsigned({reg435, (8'hb1)}))});
              reg454 = ((~|reg361) - $signed(reg443));
            end
        end
      reg455 <= $signed(reg446);
      reg456 <= {((|reg432) + {(((8'hb3) ? reg392 : wire5) * (reg439 ?
                  reg402 : wire371)),
              (~|reg439)}),
          (($signed((wire10 ^~ reg383)) || ((7'h44) ~^ (^reg444))) != (8'h9f))};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module325
#(parameter param340 = (({{(~&(7'h42)), {(8'ha4)}}} || ((((8'haf) ? (8'hac) : (8'h9d)) ? {(8'h9c)} : ((8'hb1) & (8'ha3))) ? (~((8'hbc) ? (8'hb7) : (8'hb8))) : (((8'hb9) ? (8'h9e) : (8'hb1)) ? (|(8'hbc)) : ((8'ha7) >> (8'hb6))))) > ((|(^~((8'hb0) ? (8'ha1) : (8'hac)))) ? {(((8'haa) >>> (8'hb4)) && (^~(8'hbf)))} : {{((8'hb2) ? (8'hae) : (7'h41))}, ((^(7'h44)) + (|(8'hb6)))})))
(y, clk, wire329, wire328, wire327, wire326);
  output wire [(32'h6a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire329;
  input wire [(2'h3):(1'h0)] wire328;
  input wire [(4'hf):(1'h0)] wire327;
  input wire signed [(5'h15):(1'h0)] wire326;
  wire [(5'h11):(1'h0)] wire339;
  wire [(4'ha):(1'h0)] wire338;
  wire signed [(2'h2):(1'h0)] wire337;
  wire [(4'hc):(1'h0)] wire336;
  wire signed [(4'hd):(1'h0)] wire334;
  wire [(5'h13):(1'h0)] wire333;
  wire [(5'h11):(1'h0)] wire332;
  wire signed [(3'h5):(1'h0)] wire331;
  wire signed [(3'h6):(1'h0)] wire330;
  reg [(3'h4):(1'h0)] reg335 = (1'h0);
  assign y = {wire339,
                 wire338,
                 wire337,
                 wire336,
                 wire334,
                 wire333,
                 wire332,
                 wire331,
                 wire330,
                 reg335,
                 (1'h0)};
  assign wire330 = (((($unsigned(wire326) ?
                       (wire327 * (8'hbc)) : (wire326 ?
                           wire327 : wire327)) <<< (~&{wire327})) ^~ (-wire327)) & ((^{$signed(wire327),
                       (wire329 << wire329)}) == (wire327 ?
                       (8'hb0) : $signed((8'hbe)))));
  assign wire331 = wire327[(4'h8):(2'h3)];
  assign wire332 = ($unsigned(wire331) - $unsigned(wire331));
  assign wire333 = $unsigned({{wire330}});
  assign wire334 = (^({({wire333, wire333} ?
                               $unsigned((8'ha3)) : (wire331 != wire333))} ?
                       $signed(((^~wire330) <= $unsigned(wire330))) : wire327[(4'hd):(3'h4)]));
  always
    @(posedge clk) begin
      reg335 = $unsigned($unsigned((~$signed(wire334[(4'h8):(2'h2)]))));
    end
  assign wire336 = wire330[(3'h6):(2'h2)];
  assign wire337 = wire328[(2'h3):(1'h0)];
  assign wire338 = $unsigned(wire326[(4'hc):(3'h5)]);
  assign wire339 = wire332[(4'hd):(3'h5)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module157  (y, clk, wire162, wire161, wire160, wire159, wire158);
  output wire [(32'h75d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire162;
  input wire signed [(3'h4):(1'h0)] wire161;
  input wire signed [(3'h5):(1'h0)] wire160;
  input wire [(4'hf):(1'h0)] wire159;
  input wire signed [(5'h11):(1'h0)] wire158;
  wire [(5'h10):(1'h0)] wire317;
  wire signed [(5'h10):(1'h0)] wire311;
  wire [(3'h5):(1'h0)] wire271;
  wire [(5'h10):(1'h0)] wire270;
  wire signed [(3'h6):(1'h0)] wire269;
  wire [(5'h12):(1'h0)] wire268;
  wire [(4'hc):(1'h0)] wire266;
  wire signed [(3'h5):(1'h0)] wire265;
  wire signed [(5'h10):(1'h0)] wire264;
  wire [(5'h10):(1'h0)] wire263;
  wire signed [(5'h13):(1'h0)] wire224;
  wire [(2'h2):(1'h0)] wire202;
  wire [(5'h14):(1'h0)] wire164;
  wire [(5'h13):(1'h0)] wire163;
  reg signed [(5'h13):(1'h0)] reg316 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg313 = (1'h0);
  reg signed [(4'he):(1'h0)] reg310 = (1'h0);
  reg [(4'hc):(1'h0)] reg306 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg299 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg298 = (1'h0);
  reg [(4'h9):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg296 = (1'h0);
  reg signed [(4'he):(1'h0)] reg295 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg292 = (1'h0);
  reg [(5'h11):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg286 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg283 = (1'h0);
  reg [(2'h3):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg281 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg279 = (1'h0);
  reg [(4'hb):(1'h0)] reg278 = (1'h0);
  reg [(5'h15):(1'h0)] reg275 = (1'h0);
  reg [(3'h4):(1'h0)] reg274 = (1'h0);
  reg [(5'h10):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg267 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg259 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg258 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg254 = (1'h0);
  reg [(4'h9):(1'h0)] reg252 = (1'h0);
  reg [(4'h9):(1'h0)] reg251 = (1'h0);
  reg [(5'h15):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg241 = (1'h0);
  reg [(3'h4):(1'h0)] reg240 = (1'h0);
  reg [(4'hb):(1'h0)] reg238 = (1'h0);
  reg [(2'h2):(1'h0)] reg237 = (1'h0);
  reg [(3'h5):(1'h0)] reg235 = (1'h0);
  reg [(5'h14):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg229 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg226 = (1'h0);
  reg [(2'h2):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg219 = (1'h0);
  reg [(3'h4):(1'h0)] reg214 = (1'h0);
  reg [(5'h11):(1'h0)] reg213 = (1'h0);
  reg signed [(4'he):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg207 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg200 = (1'h0);
  reg [(3'h7):(1'h0)] reg199 = (1'h0);
  reg [(5'h12):(1'h0)] reg196 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg190 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg186 = (1'h0);
  reg [(5'h14):(1'h0)] reg182 = (1'h0);
  reg [(5'h13):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg170 = (1'h0);
  reg [(3'h7):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg167 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg165 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg315 = (1'h0);
  reg [(3'h5):(1'h0)] forvar314 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar312 = (1'h0);
  reg [(4'h8):(1'h0)] reg309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg308 = (1'h0);
  reg [(4'hb):(1'h0)] forvar307 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar305 = (1'h0);
  reg signed [(4'he):(1'h0)] reg304 = (1'h0);
  reg [(4'ha):(1'h0)] forvar302 = (1'h0);
  reg [(4'hf):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg300 = (1'h0);
  reg [(4'hc):(1'h0)] forvar294 = (1'h0);
  reg [(2'h2):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar287 = (1'h0);
  reg [(4'hd):(1'h0)] reg285 = (1'h0);
  reg [(5'h11):(1'h0)] forvar284 = (1'h0);
  reg [(5'h13):(1'h0)] reg280 = (1'h0);
  reg [(4'h8):(1'h0)] forvar277 = (1'h0);
  reg [(4'hd):(1'h0)] forvar276 = (1'h0);
  reg [(4'hf):(1'h0)] reg262 = (1'h0);
  reg [(5'h13):(1'h0)] forvar261 = (1'h0);
  reg [(5'h15):(1'h0)] forvar260 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(3'h5):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar248 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg246 = (1'h0);
  reg [(4'h8):(1'h0)] reg244 = (1'h0);
  reg signed [(4'he):(1'h0)] reg243 = (1'h0);
  reg [(5'h12):(1'h0)] forvar242 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar239 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg236 = (1'h0);
  reg [(5'h14):(1'h0)] forvar233 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar227 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg222 = (1'h0);
  reg [(4'hf):(1'h0)] reg221 = (1'h0);
  reg [(5'h10):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg217 = (1'h0);
  reg [(4'h9):(1'h0)] forvar216 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar215 = (1'h0);
  reg [(3'h6):(1'h0)] reg211 = (1'h0);
  reg [(5'h15):(1'h0)] forvar210 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar206 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar204 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(5'h11):(1'h0)] reg198 = (1'h0);
  reg [(5'h13):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar194 = (1'h0);
  reg [(5'h10):(1'h0)] reg193 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg [(4'h9):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar185 = (1'h0);
  reg [(3'h4):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg181 = (1'h0);
  reg [(4'hf):(1'h0)] reg179 = (1'h0);
  reg [(4'h8):(1'h0)] forvar178 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg177 = (1'h0);
  reg [(5'h11):(1'h0)] forvar176 = (1'h0);
  reg [(4'hf):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg172 = (1'h0);
  reg [(4'hd):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar165 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar172 = (1'h0);
  reg [(4'hf):(1'h0)] reg169 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar166 = (1'h0);
  assign y = {wire317,
                 wire311,
                 wire271,
                 wire270,
                 wire269,
                 wire268,
                 wire266,
                 wire265,
                 wire264,
                 wire263,
                 wire224,
                 wire202,
                 wire164,
                 wire163,
                 reg316,
                 reg313,
                 reg310,
                 reg306,
                 reg303,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg286,
                 reg283,
                 reg282,
                 reg281,
                 reg279,
                 reg278,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg267,
                 reg259,
                 reg258,
                 reg257,
                 reg255,
                 reg254,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg247,
                 reg245,
                 reg241,
                 reg240,
                 reg238,
                 reg237,
                 reg235,
                 reg234,
                 reg232,
                 reg230,
                 reg229,
                 reg228,
                 reg226,
                 reg223,
                 reg220,
                 reg219,
                 reg214,
                 reg213,
                 reg212,
                 reg209,
                 reg208,
                 reg207,
                 reg205,
                 reg203,
                 reg200,
                 reg199,
                 reg196,
                 reg195,
                 reg190,
                 reg186,
                 reg182,
                 reg180,
                 reg174,
                 reg171,
                 reg170,
                 reg168,
                 reg167,
                 reg165,
                 reg315,
                 forvar314,
                 forvar312,
                 reg309,
                 reg308,
                 forvar307,
                 forvar305,
                 reg304,
                 forvar302,
                 reg301,
                 reg300,
                 forvar294,
                 reg289,
                 reg288,
                 forvar287,
                 reg285,
                 forvar284,
                 reg280,
                 forvar277,
                 forvar276,
                 reg262,
                 forvar261,
                 forvar260,
                 reg256,
                 reg253,
                 forvar248,
                 reg246,
                 reg244,
                 reg243,
                 forvar242,
                 forvar239,
                 reg236,
                 forvar233,
                 reg231,
                 forvar227,
                 forvar225,
                 reg222,
                 reg221,
                 reg218,
                 reg217,
                 forvar216,
                 forvar215,
                 reg211,
                 forvar210,
                 forvar206,
                 forvar204,
                 reg201,
                 reg198,
                 forvar197,
                 forvar194,
                 reg193,
                 reg192,
                 reg191,
                 reg189,
                 reg188,
                 reg187,
                 forvar185,
                 reg184,
                 reg183,
                 reg181,
                 reg179,
                 forvar178,
                 reg177,
                 forvar176,
                 reg175,
                 reg172,
                 reg166,
                 forvar165,
                 reg173,
                 forvar172,
                 reg169,
                 forvar166,
                 (1'h0)};
  assign wire163 = $signed((7'h44));
  assign wire164 = $unsigned((((wire161 ?
                           wire162[(1'h0):(1'h0)] : (wire159 && wire161)) ?
                       wire163 : {$signed(wire160),
                           (^~wire163)}) || ($unsigned(wire161[(2'h2):(1'h1)]) ?
                       {$unsigned((8'hbc)),
                           $signed(wire159)} : "spd3ecgZCOVfenCb7QTQ")));
  always
    @(posedge clk) begin
      if ((!(~^$unsigned(wire158))))
        begin
          reg165 <= (&wire162[(2'h2):(1'h0)]);
          for (forvar166 = (1'h0); (forvar166 < (2'h2)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= (8'hac);
              reg168 <= ($unsigned(wire161[(2'h3):(1'h0)]) ?
                  (forvar166[(3'h6):(3'h6)] ?
                      (((wire160 ? (8'hb6) : (8'ha0)) ?
                          (wire159 ?
                              reg165 : wire162) : ((8'ha1) != wire158)) ^ $signed(((8'hb7) ?
                          reg165 : wire160))) : "Ns0hnseumY21s8P28Aqy") : wire161);
              reg169 = ($signed({(~&wire158[(4'ha):(3'h4)])}) >= (8'hab));
              reg170 <= (reg168 >> (wire160[(2'h3):(2'h2)] && wire160));
              reg171 <= $unsigned((~({$unsigned(wire161)} ?
                  wire163[(4'h9):(1'h0)] : wire159)));
            end
          for (forvar172 = (1'h0); (forvar172 < (1'h1)); forvar172 = (forvar172 + (1'h1)))
            begin
              reg173 = reg167;
            end
        end
      else
        begin
          for (forvar165 = (1'h0); (forvar165 < (2'h3)); forvar165 = (forvar165 + (1'h1)))
            begin
              reg166 = ($signed(((-(~&reg171)) ~^ reg169)) ?
                  $unsigned($unsigned({"ESCFBF"})) : $unsigned(reg173[(4'h8):(1'h0)]));
              reg169 = "BMQQsk";
              reg170 <= ("m4L1xqz1Siy3G8" ?
                  wire164 : $signed((wire162 & wire163)));
              reg171 <= (forvar172[(4'he):(4'h9)] <<< $unsigned($signed((forvar165[(4'hc):(3'h7)] ?
                  {forvar166, forvar165} : $signed(reg168)))));
              reg172 = $signed(forvar172[(2'h3):(2'h2)]);
            end
          if ({"M",
              (wire161[(2'h2):(1'h0)] ?
                  reg173 : $signed(((wire163 ?
                      forvar172 : wire162) & ((8'hac) * (8'hac)))))})
            begin
              reg173 = ((~&(8'hba)) << $unsigned($unsigned($unsigned($unsigned(reg168)))));
              reg174 <= (({$signed((reg172 && (8'hbd)))} ?
                      wire161 : $unsigned((~|reg165))) ?
                  (~{$signed($signed(reg165)),
                      (wire160[(1'h1):(1'h1)] >= reg165[(2'h2):(1'h0)])}) : {$unsigned($unsigned((reg167 << reg168)))});
            end
          else
            begin
              reg174 <= (wire159 ?
                  (reg169[(1'h0):(1'h0)] ?
                      ((+(wire159 ? wire159 : forvar165)) ?
                          (wire164[(2'h3):(2'h2)] != reg174) : reg173[(5'h13):(4'hb)]) : (-{{wire162,
                              wire158},
                          reg168})) : (~$unsigned($unsigned({(8'hac)}))));
              reg175 = (wire159 ? (+forvar172) : (|reg168[(3'h6):(3'h4)]));
            end
          for (forvar176 = (1'h0); (forvar176 < (3'h4)); forvar176 = (forvar176 + (1'h1)))
            begin
              reg177 = "r2Mktur6SITbLrt6DCop";
            end
        end
      for (forvar178 = (1'h0); (forvar178 < (3'h4)); forvar178 = (forvar178 + (1'h1)))
        begin
          if ($signed("dCGpuzyAF"))
            begin
              reg179 = forvar178[(4'h8):(4'h8)];
              reg180 <= forvar166[(3'h6):(1'h0)];
            end
          else
            begin
              reg180 <= (8'hbc);
              reg181 = $signed({wire159});
              reg182 <= {($unsigned(({wire158, reg179} ?
                      $signed(reg174) : $unsigned((8'ha2)))) + reg175),
                  {{forvar176[(4'h9):(2'h2)]}, reg173}};
              reg183 = (-({$unsigned($signed(reg169))} ?
                  reg166[(4'hc):(2'h2)] : $signed((8'ha4))));
              reg184 = (+{wire162});
            end
          for (forvar185 = (1'h0); (forvar185 < (3'h4)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 <= {(forvar172 ?
                      ((&$unsigned(wire159)) ?
                          {forvar165,
                              reg171} : wire161) : ((^~"RpggEQARl6mVSZD5ra02") >>> {(+reg181),
                          $unsigned(reg174)}))};
            end
          reg187 = $signed(reg184[(1'h1):(1'h0)]);
          if ({$unsigned((~|$unsigned($unsigned(forvar178)))),
              (reg169 <= forvar185)})
            begin
              reg188 = $unsigned(($unsigned({reg186,
                  $signed(reg187)}) << (({forvar178,
                  (8'hbf)} + $unsigned((8'hb9))) <= reg169)));
              reg189 = ((^~(wire162 || ((wire164 ?
                  (8'ha4) : reg173) >> $signed(wire163)))) == $unsigned(($signed(wire158[(4'h8):(1'h1)]) <<< $signed(reg171[(1'h0):(1'h0)]))));
              reg190 <= ($signed((($signed(reg170) & (forvar165 ^ reg167)) >> $unsigned($unsigned(forvar165)))) - ((~(8'ha4)) <<< (8'hb0)));
              reg191 = ((~&reg190[(3'h4):(3'h4)]) ?
                  $unsigned(((^~reg183) ?
                      {(reg190 ? reg165 : wire160)} : (~{reg183,
                          (7'h40)}))) : reg179);
              reg192 = {$unsigned(($unsigned(reg184[(1'h1):(1'h1)]) ^ reg188[(3'h6):(1'h1)]))};
            end
          else
            begin
              reg190 <= $signed($signed($unsigned(forvar176[(4'he):(2'h3)])));
            end
          reg193 = reg179;
        end
      for (forvar194 = (1'h0); (forvar194 < (2'h3)); forvar194 = (forvar194 + (1'h1)))
        begin
          reg195 <= "";
          reg196 <= $signed(($unsigned(reg186[(3'h6):(1'h1)]) ?
              forvar178[(2'h3):(1'h0)] : $unsigned(reg188[(3'h4):(1'h1)])));
          for (forvar197 = (1'h0); (forvar197 < (2'h3)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 = reg179;
            end
          reg199 <= (8'hb9);
          reg200 <= (^"GhqQmIc");
        end
      reg201 = $signed((($signed(reg190[(1'h1):(1'h0)]) && (~^((8'hb4) <<< reg167))) >>> ((reg198 ?
              reg199 : (~|wire158)) ?
          ($unsigned(reg171) ?
              {forvar166, wire162} : $signed(reg187)) : (~{forvar172,
              reg179}))));
    end
  assign wire202 = (^~$unsigned({(8'h9c), (|$unsigned(reg168))}));
  always
    @(posedge clk) begin
      reg203 <= (reg167[(3'h6):(3'h6)] | (-((~&$signed((8'hbf))) ?
          ((reg165 ? wire163 : reg196) > wire202) : (~|$unsigned((8'hba))))));
      for (forvar204 = (1'h0); (forvar204 < (1'h1)); forvar204 = (forvar204 + (1'h1)))
        begin
          reg205 <= $signed({($signed((reg170 ?
                  reg180 : reg195)) >>> {$unsigned(reg195)}),
              $signed("1uVbtRCKv")});
          for (forvar206 = (1'h0); (forvar206 < (2'h2)); forvar206 = (forvar206 + (1'h1)))
            begin
              reg207 <= (^$unsigned(wire160));
              reg208 <= reg203;
            end
          reg209 <= $signed($signed($signed(wire160)));
          for (forvar210 = (1'h0); (forvar210 < (2'h3)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 = wire163;
              reg212 <= (reg190 ? reg207 : forvar210[(3'h5):(1'h1)]);
              reg213 <= (((-wire164) ?
                  (+reg167) : ($unsigned((reg211 ^~ reg174)) ?
                      ($signed(reg209) >= reg180[(4'he):(3'h4)]) : ($signed(reg196) ?
                          (~reg208) : reg186[(1'h1):(1'h1)]))) || {wire162[(3'h6):(3'h6)]});
            end
          reg214 <= ($signed($unsigned(reg205)) * $unsigned((|"aZof0yz0OTPHamE4")));
        end
      for (forvar215 = (1'h0); (forvar215 < (3'h4)); forvar215 = (forvar215 + (1'h1)))
        begin
          for (forvar216 = (1'h0); (forvar216 < (3'h4)); forvar216 = (forvar216 + (1'h1)))
            begin
              reg217 = ({reg171, $signed(wire159)} | wire162[(3'h7):(3'h7)]);
              reg218 = $signed((-(+$unsigned({reg212, reg207}))));
              reg219 <= $unsigned($signed((-"GacX8W4QYInrEe7")));
              reg220 <= ($unsigned((((^~(8'hbb)) >>> $unsigned(forvar204)) >= wire164)) < (8'ha9));
              reg221 = $signed(reg200);
            end
          reg222 = ($unsigned(reg167) ?
              $signed($unsigned(($unsigned((8'ha8)) ?
                  wire202 : (~|wire163)))) : $unsigned((^~$signed((forvar215 ?
                  reg196 : (8'h9f))))));
          reg223 <= ($unsigned((((&wire164) ?
              wire160[(2'h2):(1'h1)] : reg180) || ((^reg180) ?
              "T1SoURF4Ecltlyw" : (reg168 <= reg222)))) > {reg207[(4'hf):(4'hb)],
              reg199[(1'h0):(1'h0)]});
        end
    end
  assign wire224 = reg182[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar225 = (1'h0); (forvar225 < (1'h1)); forvar225 = (forvar225 + (1'h1)))
        begin
          reg226 <= "f7aY8L4h";
        end
      for (forvar227 = (1'h0); (forvar227 < (2'h3)); forvar227 = (forvar227 + (1'h1)))
        begin
          if ($unsigned($signed((reg174[(3'h5):(2'h3)] > (reg209[(2'h2):(1'h0)] ?
              reg219[(3'h7):(3'h5)] : reg223[(1'h0):(1'h0)])))))
            begin
              reg228 <= {(((|$signed(reg219)) < wire224[(5'h13):(4'hf)]) && (+((wire160 ?
                      (8'hb3) : wire162) <= {(8'ha2), reg226})))};
              reg229 <= $signed((+$signed(((&reg219) ?
                  (reg195 ? reg226 : wire161) : $unsigned(forvar227)))));
              reg230 <= (~|reg195);
              reg231 = (reg195[(4'h8):(2'h3)] ?
                  reg186[(1'h0):(1'h0)] : ((-((8'hb4) != reg190)) ?
                      (~|($unsigned(wire202) <<< (reg212 || (8'hba)))) : ((&(~wire160)) ^~ reg182[(5'h12):(4'he)])));
            end
          else
            begin
              reg228 <= wire160;
              reg231 = (^(-$unsigned($unsigned(wire158[(4'hc):(2'h2)]))));
              reg232 <= (!(~&$signed(reg190)));
            end
          for (forvar233 = (1'h0); (forvar233 < (3'h4)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 <= {$unsigned({reg190[(1'h0):(1'h0)]}), reg205};
              reg235 <= (reg213[(1'h1):(1'h0)] ^~ reg186);
              reg236 = $signed(forvar233[(5'h14):(5'h12)]);
            end
        end
      reg237 <= $signed(((^(((8'had) + reg229) ?
              $unsigned(reg214) : {wire158, (8'hb6)})) ?
          $signed((~&$unsigned((8'hae)))) : (~^(8'hb6))));
      reg238 <= (|(~^(wire160[(3'h4):(2'h2)] > reg220[(1'h0):(1'h0)])));
      for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
        begin
          reg240 <= reg207[(4'hd):(3'h4)];
          reg241 <= $signed("DE2fHM6KlSD8JIAIMOL");
          for (forvar242 = (1'h0); (forvar242 < (1'h0)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 = reg195;
              reg244 = {(wire161[(2'h2):(1'h1)] ?
                      reg231[(1'h0):(1'h0)] : reg190[(3'h6):(3'h4)])};
              reg245 <= ((~^(^($unsigned((7'h42)) ?
                  (wire159 * reg240) : reg244))) ^~ {(~&$signed((wire224 - reg237)))});
              reg246 = {reg230[(3'h6):(2'h2)]};
              reg247 <= (($signed(({wire159} > reg167)) * ($signed((forvar233 ?
                  wire163 : (8'hb4))) + (~^{reg214,
                  reg243}))) ^ reg226[(3'h7):(3'h4)]);
            end
          for (forvar248 = (1'h0); (forvar248 < (2'h2)); forvar248 = (forvar248 + (1'h1)))
            begin
              reg249 <= $unsigned((-$signed($unsigned($signed(reg231)))));
              reg250 <= reg236[(3'h7):(3'h4)];
              reg251 <= ($unsigned((((reg245 ?
                          reg229 : reg226) >= $signed(reg205)) ?
                      (((8'ha7) >= reg196) && (|reg244)) : $signed($unsigned(wire162)))) ?
                  "IJnHLPfKIiF" : $signed({(|{(8'hbc)}), ""}));
              reg252 <= reg186[(1'h1):(1'h0)];
              reg253 = reg182;
            end
          if ({$unsigned(forvar239)})
            begin
              reg254 <= ("lDNFNYFv9zGN" ?
                  $signed(reg199) : (reg209[(2'h3):(2'h3)] || reg208[(4'he):(3'h4)]));
              reg255 <= ($unsigned((|(reg252 << (forvar233 ?
                  wire161 : reg238)))) > $signed(wire202));
            end
          else
            begin
              reg254 <= reg199[(3'h4):(1'h1)];
              reg256 = (8'hb0);
              reg257 <= forvar248;
              reg258 <= $signed($unsigned(reg257));
            end
        end
    end
  always
    @(posedge clk) begin
      reg259 <= "M790cOCZ527UJqB";
      for (forvar260 = (1'h0); (forvar260 < (1'h1)); forvar260 = (forvar260 + (1'h1)))
        begin
          for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
            begin
              reg262 = $signed(forvar260[(5'h15):(4'hf)]);
            end
        end
    end
  assign wire263 = $unsigned(({(wire162 ?
                           reg167[(3'h4):(1'h1)] : $signed(reg250))} >= ((((8'hbb) ?
                           reg165 : reg247) && wire159) ?
                       "" : reg165)));
  assign wire264 = {$unsigned(wire160)};
  assign wire265 = $unsigned(wire164[(3'h7):(1'h0)]);
  assign wire266 = {(reg212 ?
                           {$unsigned($unsigned(reg171))} : $unsigned(reg182)),
                       reg223};
  always
    @(posedge clk) begin
      reg267 <= (reg251 ^ $signed({"T"}));
    end
  assign wire268 = wire161[(2'h3):(2'h3)];
  assign wire269 = $unsigned(($signed(reg171) >= ((wire266 ?
                       (reg205 << wire164) : wire265) >= reg212)));
  assign wire270 = "sQ3Jkvg8QxU4BGt";
  assign wire271 = reg229[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      reg272 <= reg171[(2'h3):(2'h3)];
      reg273 <= (8'ha6);
      reg274 <= wire161[(2'h2):(2'h2)];
      reg275 <= $signed({reg273, reg255});
    end
  always
    @(posedge clk) begin
      for (forvar276 = (1'h0); (forvar276 < (2'h3)); forvar276 = (forvar276 + (1'h1)))
        begin
          for (forvar277 = (1'h0); (forvar277 < (2'h3)); forvar277 = (forvar277 + (1'h1)))
            begin
              reg278 <= wire263;
              reg279 <= (reg250[(5'h15):(4'he)] & (reg235 ?
                  wire162 : $unsigned($signed($signed(wire271)))));
            end
          if (((^~reg207[(4'ha):(4'h9)]) ?
              (^~{((reg186 ? (8'ha6) : reg186) | reg274),
                  ((8'ha0) ? reg219 : (reg247 ? reg167 : reg226))}) : reg212))
            begin
              reg280 = (^~(reg279[(1'h1):(1'h1)] ?
                  (forvar276 ?
                      ((reg279 ? reg186 : (8'h9c)) ?
                          (-forvar277) : wire224[(4'ha):(4'ha)]) : "T1u") : wire159[(2'h3):(1'h1)]));
              reg281 <= (wire268 ?
                  $unsigned(reg207[(1'h1):(1'h1)]) : (reg235[(1'h1):(1'h1)] ?
                      (^(forvar276 ? reg228 : reg165)) : ($signed((wire266 ?
                          reg223 : forvar277)) * ((reg205 < reg241) ?
                          reg170[(4'ha):(3'h4)] : $signed(wire266)))));
              reg282 <= {$unsigned(reg168)};
            end
          else
            begin
              reg280 = (~(reg252 ? reg273 : reg238[(1'h0):(1'h0)]));
              reg281 <= ({wire271} ?
                  $unsigned((wire224[(3'h4):(3'h4)] ?
                      ($signed((7'h42)) - "3NfXZXu3uZyQJp") : $signed((8'ha7)))) : ((reg200[(3'h4):(3'h4)] ?
                      $signed((|reg229)) : (|$unsigned(forvar277))) != ({forvar277} ?
                      reg186[(3'h7):(1'h1)] : (wire202 ?
                          (~|reg232) : (-reg258)))));
              reg282 <= "lXy4KqW0r0z";
            end
          reg283 <= $signed({"33kM"});
          for (forvar284 = (1'h0); (forvar284 < (1'h0)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 = reg258;
              reg286 <= reg249[(5'h10):(4'ha)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar287 = (1'h0); (forvar287 < (3'h4)); forvar287 = (forvar287 + (1'h1)))
        begin
          if ($signed({(reg219 ? reg257 : wire164),
              (reg180 - {$signed(wire164)})}))
            begin
              reg288 = (~^(^(8'ha4)));
              reg289 = reg213;
              reg290 <= reg288[(4'ha):(1'h0)];
              reg291 <= $signed((8'hb1));
            end
          else
            begin
              reg290 <= {(wire158 >> $unsigned(reg214))};
              reg291 <= ((|(~&"WXzrt6T7FF")) <= (((^~$signed(reg240)) >>> reg207[(1'h1):(1'h0)]) == $signed(((reg196 ?
                      reg174 : reg219) ?
                  reg182[(4'ha):(3'h4)] : (~&reg273)))));
              reg292 <= ((8'haa) ?
                  wire265[(1'h0):(1'h0)] : (({(8'ha4)} ?
                      reg190 : $unsigned({(8'hba),
                          reg278})) == $unsigned(reg289)));
            end
          reg293 <= reg212;
          for (forvar294 = (1'h0); (forvar294 < (1'h0)); forvar294 = (forvar294 + (1'h1)))
            begin
              reg295 <= (wire158[(1'h1):(1'h0)] <= ($signed($unsigned($signed((8'ha4)))) ?
                  (-{(&wire159),
                      $signed(reg209)}) : $signed(({reg190} < (reg275 * reg245)))));
              reg296 <= $signed($unsigned(((|(~^reg182)) ?
                  (wire159[(4'he):(4'h8)] ?
                      (wire164 ?
                          wire202 : reg170) : {reg241}) : (~&$signed(reg196)))));
            end
          if ($unsigned(($unsigned(((+reg292) ?
              (~&wire162) : ((8'h9c) == reg226))) ~^ (+$signed($unsigned(reg289))))))
            begin
              reg297 <= (reg240 - (reg249 > ($signed(reg250[(3'h5):(1'h0)]) ?
                  {(reg257 <= reg208),
                      $unsigned(reg267)} : "R0gEWxA9AfLxBEU2GNq")));
            end
          else
            begin
              reg297 <= (((((wire163 <= reg234) ~^ reg297) & (^~(!wire163))) || $signed($signed($unsigned(reg282)))) ?
                  wire265 : reg254);
              reg298 <= reg245;
            end
        end
      if ("xRzOLGgTYs31UlwZu4")
        begin
          reg299 <= $signed("oI7sePO0IIJi");
          reg300 = wire161[(1'h0):(1'h0)];
        end
      else
        begin
          if (reg288)
            begin
              reg300 = reg289[(2'h2):(1'h1)];
              reg301 = {($signed((((8'hbe) && reg171) ?
                      $unsigned(reg168) : (&reg282))) <= $unsigned(reg223)),
                  reg223[(1'h1):(1'h1)]};
            end
          else
            begin
              reg300 = $unsigned((reg240 != reg300[(2'h3):(1'h0)]));
              reg301 = reg168[(3'h7):(3'h7)];
            end
          for (forvar302 = (1'h0); (forvar302 < (3'h4)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg303 <= $unsigned((~&$unsigned($signed({(8'hbd), (8'ha4)}))));
            end
          reg304 = reg258;
        end
      for (forvar305 = (1'h0); (forvar305 < (2'h3)); forvar305 = (forvar305 + (1'h1)))
        begin
          reg306 <= (~(|((reg245 ?
                  $unsigned(reg195) : (reg232 ? reg273 : (8'ha3))) ?
              (+(~|wire271)) : $unsigned((reg286 ? (8'hbd) : reg252)))));
          for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
            begin
              reg308 = (+$signed("pYq0RrBQW6u6"));
              reg309 = (~&$signed($unsigned(({reg168, (8'hb2)} & (~|reg255)))));
            end
          reg310 <= "l";
        end
    end
  assign wire311 = $unsigned(($signed($signed((reg214 ^ reg174))) || $unsigned((~&reg299))));
  always
    @(posedge clk) begin
      for (forvar312 = (1'h0); (forvar312 < (3'h4)); forvar312 = (forvar312 + (1'h1)))
        begin
          reg313 <= $signed(reg259[(1'h0):(1'h0)]);
        end
      for (forvar314 = (1'h0); (forvar314 < (2'h2)); forvar314 = (forvar314 + (1'h1)))
        begin
          if ((8'hb7))
            begin
              reg315 = (((|(reg195 ?
                      (reg278 ?
                          reg208 : reg310) : reg186[(1'h0):(1'h0)])) >= wire162[(1'h0):(1'h0)]) ?
                  $unsigned(reg259) : reg257);
            end
          else
            begin
              reg316 <= (~&(-($unsigned(reg255) << reg232)));
            end
        end
    end
  assign wire317 = (wire163[(3'h5):(3'h4)] ?
                       $signed((reg247 ?
                           $unsigned((reg237 >>> reg229)) : $unsigned((reg241 ?
                               (8'hbf) : reg273)))) : ({$unsigned(reg199[(3'h5):(2'h3)]),
                               $unsigned((wire161 ? reg258 : (8'hb2)))} ?
                           reg306[(3'h6):(3'h4)] : reg257));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module134  (y, clk, wire139, wire138, wire137, wire136, wire135);
  output wire [(32'h77):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire139;
  input wire [(2'h3):(1'h0)] wire138;
  input wire signed [(4'he):(1'h0)] wire137;
  input wire signed [(5'h11):(1'h0)] wire136;
  input wire [(4'hd):(1'h0)] wire135;
  wire [(3'h6):(1'h0)] wire150;
  wire signed [(5'h13):(1'h0)] wire149;
  wire [(5'h12):(1'h0)] wire148;
  wire signed [(4'h9):(1'h0)] wire147;
  reg [(3'h5):(1'h0)] reg145 = (1'h0);
  reg [(2'h3):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg142 = (1'h0);
  reg [(4'h8):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg143 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar141 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar140 = (1'h0);
  assign y = {wire150,
                 wire149,
                 wire148,
                 wire147,
                 reg145,
                 reg144,
                 reg142,
                 reg146,
                 reg143,
                 forvar141,
                 forvar140,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar140 = (1'h0); (forvar140 < (3'h4)); forvar140 = (forvar140 + (1'h1)))
        begin
          for (forvar141 = (1'h0); (forvar141 < (2'h2)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg142 <= ((+($signed(forvar141) + ((~&forvar140) < (wire135 ^ wire139)))) ?
                  (wire137 ?
                      ($signed(wire137[(4'hd):(1'h1)]) != $unsigned($signed((8'hba)))) : ($signed({forvar140}) >>> $unsigned((^~wire136)))) : forvar141[(1'h0):(1'h0)]);
              reg143 = $signed(reg142);
              reg144 <= reg142[(3'h4):(1'h1)];
              reg145 <= reg142[(2'h2):(1'h0)];
            end
          reg146 = reg144;
        end
    end
  assign wire147 = (&$signed($signed(reg145[(3'h4):(2'h2)])));
  assign wire148 = {{wire138[(1'h1):(1'h0)], (!$signed($signed(wire135)))}};
  assign wire149 = (~|$unsigned($signed(reg145)));
  assign wire150 = (^~{(~^((wire149 ? (8'ha6) : reg142) <<< (~^reg144)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module11
#(parameter param129 = (^~(((8'hb5) - (^~((8'hb2) ? (8'hab) : (8'haf)))) ? (^(7'h44)) : {(+(~&(8'haa)))})), 
parameter param130 = param129)
(y, clk, wire16, wire15, wire14, wire13, wire12);
  output wire [(32'h540):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire16;
  input wire signed [(4'hd):(1'h0)] wire15;
  input wire signed [(3'h5):(1'h0)] wire14;
  input wire [(5'h12):(1'h0)] wire13;
  input wire [(4'hf):(1'h0)] wire12;
  wire [(4'h9):(1'h0)] wire128;
  wire signed [(5'h14):(1'h0)] wire69;
  wire signed [(4'hf):(1'h0)] wire68;
  wire [(4'h9):(1'h0)] wire67;
  wire signed [(3'h4):(1'h0)] wire66;
  wire signed [(5'h15):(1'h0)] wire18;
  wire signed [(2'h3):(1'h0)] wire17;
  reg [(3'h7):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg124 = (1'h0);
  reg [(5'h14):(1'h0)] reg123 = (1'h0);
  reg [(4'h9):(1'h0)] reg121 = (1'h0);
  reg [(5'h14):(1'h0)] reg120 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg [(4'hd):(1'h0)] reg117 = (1'h0);
  reg [(5'h10):(1'h0)] reg115 = (1'h0);
  reg [(5'h15):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  reg [(4'h8):(1'h0)] reg112 = (1'h0);
  reg [(3'h6):(1'h0)] reg110 = (1'h0);
  reg [(5'h10):(1'h0)] reg107 = (1'h0);
  reg [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg102 = (1'h0);
  reg [(5'h13):(1'h0)] reg99 = (1'h0);
  reg [(3'h7):(1'h0)] reg97 = (1'h0);
  reg [(4'h9):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg94 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg91 = (1'h0);
  reg [(4'hf):(1'h0)] reg90 = (1'h0);
  reg [(4'hd):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg87 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg86 = (1'h0);
  reg [(4'hd):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg84 = (1'h0);
  reg [(4'hc):(1'h0)] reg82 = (1'h0);
  reg [(3'h7):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(3'h7):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg63 = (1'h0);
  reg [(2'h2):(1'h0)] reg60 = (1'h0);
  reg [(5'h11):(1'h0)] reg59 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg55 = (1'h0);
  reg [(5'h12):(1'h0)] reg54 = (1'h0);
  reg [(3'h6):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg52 = (1'h0);
  reg signed [(4'he):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg50 = (1'h0);
  reg [(5'h13):(1'h0)] reg49 = (1'h0);
  reg [(3'h7):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg38 = (1'h0);
  reg [(2'h3):(1'h0)] reg46 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg44 = (1'h0);
  reg [(5'h12):(1'h0)] reg43 = (1'h0);
  reg signed [(4'he):(1'h0)] reg42 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg39 = (1'h0);
  reg [(5'h15):(1'h0)] reg35 = (1'h0);
  reg [(2'h3):(1'h0)] reg34 = (1'h0);
  reg [(4'ha):(1'h0)] reg28 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg27 = (1'h0);
  reg [(5'h12):(1'h0)] reg25 = (1'h0);
  reg [(4'ha):(1'h0)] reg24 = (1'h0);
  reg [(4'hf):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg22 = (1'h0);
  reg [(5'h10):(1'h0)] reg21 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar125 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg116 = (1'h0);
  reg [(2'h3):(1'h0)] forvar111 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar109 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar108 = (1'h0);
  reg [(5'h14):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg104 = (1'h0);
  reg [(5'h11):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg101 = (1'h0);
  reg [(3'h7):(1'h0)] forvar100 = (1'h0);
  reg [(4'hf):(1'h0)] reg98 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar93 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg92 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar83 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar78 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar77 = (1'h0);
  reg [(4'hd):(1'h0)] reg74 = (1'h0);
  reg [(4'h8):(1'h0)] reg73 = (1'h0);
  reg [(3'h6):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar71 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar70 = (1'h0);
  reg [(4'he):(1'h0)] reg62 = (1'h0);
  reg [(5'h15):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg57 = (1'h0);
  reg [(5'h12):(1'h0)] forvar56 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg45 = (1'h0);
  reg [(3'h4):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar38 = (1'h0);
  reg [(4'h9):(1'h0)] reg37 = (1'h0);
  reg [(5'h14):(1'h0)] forvar36 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg33 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg30 = (1'h0);
  reg [(4'hb):(1'h0)] forvar29 = (1'h0);
  reg [(5'h11):(1'h0)] forvar26 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar20 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar19 = (1'h0);
  assign y = {wire128,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire18,
                 wire17,
                 reg126,
                 reg124,
                 reg123,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg110,
                 reg107,
                 reg106,
                 reg103,
                 reg102,
                 reg99,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg91,
                 reg90,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg76,
                 reg75,
                 reg65,
                 reg64,
                 reg63,
                 reg60,
                 reg59,
                 reg58,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg38,
                 reg46,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg39,
                 reg35,
                 reg34,
                 reg28,
                 reg27,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg127,
                 forvar125,
                 reg122,
                 reg116,
                 forvar111,
                 forvar109,
                 forvar108,
                 reg105,
                 reg104,
                 reg93,
                 reg101,
                 forvar100,
                 reg98,
                 forvar93,
                 reg92,
                 reg89,
                 forvar83,
                 forvar78,
                 forvar77,
                 reg74,
                 reg73,
                 reg72,
                 forvar71,
                 forvar70,
                 reg62,
                 reg61,
                 reg57,
                 forvar56,
                 reg45,
                 reg40,
                 forvar38,
                 reg37,
                 forvar36,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 forvar26,
                 forvar20,
                 forvar19,
                 (1'h0)};
  assign wire17 = (wire15[(1'h1):(1'h1)] ?
                      $unsigned($signed($signed("lqNfo"))) : wire16[(4'hf):(3'h6)]);
  assign wire18 = $unsigned($signed($signed(({wire12} ?
                      $unsigned(wire15) : wire12))));
  always
    @(posedge clk) begin
      for (forvar19 = (1'h0); (forvar19 < (1'h0)); forvar19 = (forvar19 + (1'h1)))
        begin
          for (forvar20 = (1'h0); (forvar20 < (1'h1)); forvar20 = (forvar20 + (1'h1)))
            begin
              reg21 <= $unsigned({$unsigned(wire15)});
              reg22 <= forvar19[(2'h3):(2'h2)];
              reg23 <= $signed(wire14);
              reg24 <= (|wire18[(5'h14):(4'hd)]);
            end
        end
      reg25 <= $signed((~$unsigned((^$unsigned(wire14)))));
      for (forvar26 = (1'h0); (forvar26 < (3'h4)); forvar26 = (forvar26 + (1'h1)))
        begin
          reg27 <= (((wire12[(2'h2):(1'h0)] < ((reg24 ?
                  wire18 : (8'had)) ^~ (reg22 == wire12))) ?
              $unsigned((~^(wire16 == (8'had)))) : (-$signed((~|reg23)))) >> $signed(reg23[(3'h5):(1'h0)]));
          reg28 <= ({reg22, (8'ha4)} ?
              ($signed(reg27) ?
                  (~&$signed($unsigned(wire16))) : ($signed((8'hb0)) >= ((reg25 ?
                      reg25 : wire12) ^ (wire18 & reg27)))) : ($unsigned($unsigned($signed((7'h44)))) ?
                  $signed(wire17[(1'h0):(1'h0)]) : $signed(((reg23 ?
                      (8'hbd) : wire18) - (8'hbe)))));
          for (forvar29 = (1'h0); (forvar29 < (1'h1)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 = (($signed($unsigned({wire12})) > $signed(reg24[(1'h0):(1'h0)])) ?
                  ("v33aAeXRP1W" < reg24[(1'h1):(1'h1)]) : ({reg24,
                      forvar20[(5'h13):(4'he)]} - $signed(reg23)));
              reg31 = (~$unsigned($unsigned(((wire18 || reg23) ?
                  (~|reg28) : reg24[(3'h4):(1'h1)]))));
            end
          reg32 = ((forvar29 || wire14[(2'h3):(2'h3)]) ?
              $signed($signed({wire15})) : wire12[(4'h8):(3'h7)]);
        end
    end
  always
    @(posedge clk) begin
      reg33 = $unsigned($unsigned((~|$signed((wire18 || wire13)))));
      reg34 <= ((|reg23[(4'hf):(4'ha)]) ?
          (8'h9c) : (wire12 << ($signed(wire14) ?
              (wire15 ?
                  reg25 : (7'h41)) : (wire13[(1'h0):(1'h0)] | (^~reg22)))));
      reg35 <= wire17[(1'h1):(1'h1)];
      if ($unsigned((7'h41)))
        begin
          for (forvar36 = (1'h0); (forvar36 < (2'h3)); forvar36 = (forvar36 + (1'h1)))
            begin
              reg37 = reg33;
            end
          for (forvar38 = (1'h0); (forvar38 < (1'h1)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= ({(&$unsigned({reg21}))} ?
                  reg28 : (-($signed(reg22[(2'h3):(1'h1)]) == {(wire17 <= (8'ha8))})));
              reg40 = wire15[(3'h7):(3'h4)];
              reg41 <= (wire15 <= wire12);
            end
          reg42 <= ((!"IDKTmkD") & (8'ha1));
          if ({forvar36})
            begin
              reg43 <= $unsigned($unsigned($signed((|(reg37 <= wire15)))));
            end
          else
            begin
              reg43 <= $unsigned(reg27);
              reg44 <= {$signed(reg43[(3'h6):(2'h3)])};
              reg45 = ($unsigned(wire18[(1'h0):(1'h0)]) <= wire17);
              reg46 <= (^~$signed((&$signed(reg21))));
            end
        end
      else
        begin
          for (forvar36 = (1'h0); (forvar36 < (3'h4)); forvar36 = (forvar36 + (1'h1)))
            begin
              reg38 <= wire12[(4'hc):(3'h7)];
              reg40 = ($signed($signed((^~reg33[(3'h6):(2'h3)]))) + $unsigned(reg42[(2'h2):(2'h2)]));
              reg41 <= $signed((reg39 && (($signed((8'ha5)) ?
                      wire12[(4'hc):(4'hc)] : $signed(reg38)) ?
                  (^~$unsigned(reg41)) : wire14)));
              reg42 <= $signed(reg25);
              reg43 <= (8'ha5);
            end
          if ($signed($unsigned(reg38[(4'he):(2'h2)])))
            begin
              reg45 = (reg27[(3'h4):(1'h1)] ?
                  "66BkN55qDXaRD" : (wire18[(5'h12):(2'h3)] ?
                      $signed(((forvar38 ? forvar36 : reg42) > (reg44 ?
                          reg38 : wire13))) : $signed(($unsigned(wire15) ?
                          $unsigned((8'hb6)) : $unsigned(reg46)))));
              reg46 <= ((~&$signed((~&(|reg27)))) ?
                  (({"sOSJ7h", (~^(8'hae))} - {reg42}) < (((8'ha8) ?
                          reg35 : $unsigned(wire17)) ?
                      (((8'hb7) ? (8'ha8) : wire14) != (reg25 ?
                          reg28 : wire16)) : $unsigned((reg28 < (8'ha6))))) : {reg39});
              reg47 <= $unsigned(reg44[(2'h3):(2'h2)]);
              reg48 <= reg21[(4'hf):(1'h0)];
            end
          else
            begin
              reg44 <= $unsigned(({$unsigned(wire13)} ?
                  $signed($signed($signed(reg47))) : ({forvar38[(3'h7):(2'h3)],
                      (reg21 || reg28)} <= {$unsigned(forvar36),
                      (reg42 && wire18)})));
              reg46 <= ($signed(wire14[(3'h4):(3'h4)]) << $unsigned(reg40[(2'h3):(2'h2)]));
              reg47 <= ((|(~^{wire14[(3'h5):(3'h4)]})) ?
                  ((^~$signed($signed(reg42))) ?
                      (($signed((8'h9e)) - (reg39 ? wire18 : reg47)) ?
                          $signed((reg40 ?
                              forvar38 : reg42)) : reg43[(1'h0):(1'h0)]) : {(+$signed(reg25))}) : $unsigned(reg44[(2'h2):(2'h2)]));
              reg48 <= "38gtf";
              reg49 <= $unsigned(($signed(wire18) <= $signed($unsigned((reg43 ^~ reg44)))));
            end
          reg50 <= (|((wire13 ? (wire17 > (~reg42)) : (!$unsigned(reg40))) ?
              wire18 : forvar36));
          if ($signed($unsigned($signed(((reg43 ? reg21 : forvar38) ?
              reg48[(1'h1):(1'h1)] : (reg22 != forvar38))))))
            begin
              reg51 <= reg40;
              reg52 <= (wire16[(2'h2):(2'h2)] >= $signed($signed(wire16)));
            end
          else
            begin
              reg51 <= {(~|$signed($signed((wire14 > reg41)))),
                  {($unsigned($signed(reg33)) && reg27[(2'h3):(1'h1)])}};
              reg52 <= $unsigned({($unsigned((+wire14)) ?
                      reg21 : $signed($signed(wire12))),
                  (8'hb3)});
              reg53 <= (~^(~&wire12));
              reg54 <= wire16;
            end
          reg55 <= $unsigned($unsigned((~|($unsigned(reg49) && wire17))));
        end
      for (forvar56 = (1'h0); (forvar56 < (1'h1)); forvar56 = (forvar56 + (1'h1)))
        begin
          reg57 = reg47[(2'h3):(2'h3)];
          if (forvar36)
            begin
              reg58 <= wire18[(4'hb):(2'h2)];
              reg59 <= $signed((7'h40));
              reg60 <= $unsigned((&((~^{wire17}) ?
                  $signed(reg39[(1'h1):(1'h0)]) : $signed(reg42))));
              reg61 = (~|(($unsigned(reg37[(3'h6):(3'h5)]) ?
                      (~(reg41 ^ wire16)) : forvar56[(3'h6):(3'h5)]) ?
                  {$unsigned((8'ha3)),
                      ((reg55 + wire16) + (8'h9c))} : ($unsigned((^reg59)) == ($signed(reg53) ?
                      reg60[(2'h2):(2'h2)] : forvar36[(3'h6):(2'h3)]))));
              reg62 = reg25[(3'h7):(2'h3)];
            end
          else
            begin
              reg61 = {$signed($unsigned(("X4YzRodclRG" != ((8'ha0) < reg48)))),
                  forvar56};
              reg63 <= (~(reg48 ?
                  {$unsigned($signed(forvar36))} : reg42[(4'hc):(2'h3)]));
            end
          reg64 <= $signed(reg24);
        end
    end
  always
    @(posedge clk) begin
      reg65 <= reg51[(3'h7):(2'h3)];
    end
  assign wire66 = {(~&{$unsigned((|reg41))})};
  assign wire67 = ((8'ha4) ?
                      ((^((reg58 | reg34) & ((8'h9d) ^ reg41))) > wire14[(2'h3):(2'h2)]) : reg43);
  assign wire68 = ($unsigned((^{reg63[(4'h8):(3'h4)], $unsigned(reg52)})) ?
                      (^~(^{(wire12 - reg51)})) : (!wire66[(3'h4):(1'h1)]));
  assign wire69 = (8'ha5);
  always
    @(posedge clk) begin
      for (forvar70 = (1'h0); (forvar70 < (2'h3)); forvar70 = (forvar70 + (1'h1)))
        begin
          for (forvar71 = (1'h0); (forvar71 < (3'h4)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 = (($unsigned(wire69[(3'h7):(1'h1)]) ^ ({(reg60 <= reg28),
                          $unsigned(reg24)} ?
                      $signed((reg25 ? (8'had) : reg53)) : (^(reg53 ?
                          wire13 : wire18)))) ?
                  wire15[(1'h1):(1'h0)] : $signed($unsigned(wire12)));
              reg73 = reg65[(4'hc):(2'h3)];
              reg74 = ((!$unsigned((~^wire68[(4'hb):(3'h6)]))) ^ ($signed((~(reg50 == wire12))) && $unsigned("e0YFTR0ikaLx7gVs89Oy")));
              reg75 <= $signed($unsigned(reg27));
              reg76 <= ($unsigned((~($unsigned(reg51) ? {forvar71} : reg21))) ?
                  (!(reg73 >= $unsigned($signed((7'h44))))) : ((-reg47) ?
                      ($signed($signed(reg58)) ~^ wire13[(1'h1):(1'h0)]) : reg74));
            end
        end
      for (forvar77 = (1'h0); (forvar77 < (3'h4)); forvar77 = (forvar77 + (1'h1)))
        begin
          for (forvar78 = (1'h0); (forvar78 < (2'h2)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 <= ((~|$signed($signed(reg28[(3'h4):(3'h4)]))) ?
                  $unsigned("Wt4Lp1") : ($unsigned(($unsigned(reg44) ?
                          $signed(reg48) : {wire15, (8'hbc)})) ?
                      (!(!(reg41 ? reg52 : wire16))) : ((~&$signed(reg55)) ?
                          (&$signed(reg25)) : $unsigned((~&reg60)))));
            end
          reg80 <= wire15[(2'h3):(1'h0)];
          reg81 <= $unsigned(reg49[(4'h9):(4'h8)]);
          reg82 <= (|wire16[(1'h1):(1'h1)]);
        end
      for (forvar83 = (1'h0); (forvar83 < (2'h3)); forvar83 = (forvar83 + (1'h1)))
        begin
          reg84 <= $unsigned(reg51);
          if ((8'had))
            begin
              reg85 <= (((^($unsigned(wire16) ? (|(8'ha5)) : (~&reg82))) ?
                  $unsigned(reg73[(4'h8):(1'h0)]) : (~reg81[(3'h7):(2'h2)])) & $unsigned(reg47));
              reg86 <= $unsigned({{((~wire17) ~^ reg34), reg82},
                  (({reg44} <<< reg44) ? (8'hae) : wire66[(3'h4):(2'h3)])});
            end
          else
            begin
              reg85 <= $unsigned({$unsigned((~&(reg51 ? wire66 : forvar83)))});
            end
          if ($unsigned(forvar78[(3'h5):(2'h3)]))
            begin
              reg87 <= $signed(reg85);
              reg88 <= {reg75[(2'h2):(1'h0)], reg82[(2'h2):(2'h2)]};
            end
          else
            begin
              reg89 = wire16[(2'h3):(2'h2)];
              reg90 <= {(wire69[(1'h1):(1'h1)] <= $unsigned($unsigned((reg89 ?
                      forvar77 : (8'haa)))))};
            end
          reg91 <= reg39[(2'h2):(2'h2)];
          reg92 = (|$unsigned((wire18 * ((reg89 <<< (8'haa)) ?
              (forvar77 ? reg63 : reg88) : (|reg25)))));
        end
      if ($signed(wire66[(2'h3):(2'h2)]))
        begin
          for (forvar93 = (1'h0); (forvar93 < (1'h0)); forvar93 = (forvar93 + (1'h1)))
            begin
              reg94 <= $signed(reg44);
              reg95 <= reg49;
            end
          reg96 <= $unsigned($signed($unsigned((~^$signed(reg55)))));
          if ((~|(~&reg89)))
            begin
              reg97 <= forvar83;
              reg98 = ((8'hb2) ?
                  ((((reg90 ?
                          reg44 : (8'hba)) ~^ (|reg86)) * $unsigned($signed(reg87))) ?
                      {(~$unsigned(reg87))} : reg92[(1'h0):(1'h0)]) : (8'ha7));
            end
          else
            begin
              reg97 <= wire14;
              reg99 <= ($signed((({(8'had)} ?
                          (reg51 ? reg76 : (8'hb6)) : $unsigned(wire67)) ?
                      reg50 : $signed($signed(reg81)))) ?
                  (8'hbf) : (-$signed(reg28)));
            end
          for (forvar100 = (1'h0); (forvar100 < (2'h3)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 = $unsigned($unsigned($signed({(reg86 >> forvar78),
                  $signed(reg24)})));
              reg102 <= $unsigned((~|$unsigned({(~^(8'haf)), {reg73, reg58}})));
            end
          reg103 <= reg54[(5'h11):(4'ha)];
        end
      else
        begin
          reg93 = $unsigned($unsigned(($unsigned(reg50) < $signed(reg103[(2'h3):(1'h0)]))));
          reg98 = $unsigned({({(reg34 & reg47),
                  reg60[(2'h2):(1'h1)]} < $unsigned(reg34[(2'h2):(1'h0)])),
              reg88});
          reg99 <= $signed((7'h41));
          for (forvar100 = (1'h0); (forvar100 < (2'h2)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 = reg96;
              reg104 = reg75[(2'h3):(2'h3)];
              reg105 = reg103[(3'h7):(2'h2)];
              reg106 <= reg73[(3'h7):(3'h7)];
            end
          reg107 <= (|((8'ha3) ?
              ((~|(~reg28)) < $signed((reg41 ?
                  (8'hb4) : (8'h9f)))) : forvar78[(1'h0):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      for (forvar108 = (1'h0); (forvar108 < (2'h2)); forvar108 = (forvar108 + (1'h1)))
        begin
          for (forvar109 = (1'h0); (forvar109 < (2'h2)); forvar109 = (forvar109 + (1'h1)))
            begin
              reg110 <= $unsigned($signed((8'had)));
            end
          for (forvar111 = (1'h0); (forvar111 < (2'h2)); forvar111 = (forvar111 + (1'h1)))
            begin
              reg112 <= ((wire67[(1'h0):(1'h0)] ?
                  {$signed($signed(reg82)),
                      ($unsigned(reg42) * {reg90})} : (~&reg27[(1'h1):(1'h0)])) + ({(reg85 && (reg64 ?
                      reg21 : reg110))} ~^ ($unsigned({(8'ha6),
                  reg80}) & reg91)));
              reg113 <= reg34;
              reg114 <= {wire12};
            end
          if ((~&$unsigned($signed((wire12[(4'hb):(3'h7)] ?
              (reg47 ? reg43 : reg64) : reg88)))))
            begin
              reg115 <= $unsigned({reg86});
              reg116 = ({reg42,
                  ((^(reg27 << reg114)) ?
                      (reg35 ?
                          reg115 : $signed(reg65)) : $signed($signed(wire15)))} ^~ reg41);
              reg117 <= "dufOmeBfxSuZgq";
            end
          else
            begin
              reg115 <= forvar109[(2'h3):(2'h3)];
              reg117 <= (reg63 ?
                  ($unsigned(((wire15 * (8'hb6)) ^ $unsigned(reg102))) ?
                      $unsigned((reg35[(4'hc):(3'h6)] ?
                          (8'h9c) : wire69)) : (~(reg114[(3'h6):(3'h5)] != (reg59 & reg41)))) : "KoRUxX3Z9");
              reg118 <= (~^reg22[(2'h3):(1'h1)]);
              reg119 <= reg51[(3'h6):(1'h1)];
              reg120 <= wire13;
            end
          reg121 <= reg34[(2'h3):(1'h1)];
          reg122 = {reg76[(2'h3):(1'h0)],
              (({reg24[(4'h8):(3'h4)],
                      forvar108} - $signed(reg54[(4'he):(2'h2)])) ?
                  ((8'hb0) ?
                      $unsigned(wire16[(5'h10):(4'h9)]) : ((|(8'hb9)) ?
                          wire68 : reg106)) : reg50)};
        end
      reg123 <= (&$signed(reg44[(1'h0):(1'h0)]));
      reg124 <= (+(reg115[(4'hc):(1'h1)] ?
          $signed($unsigned((^reg47))) : {reg44[(2'h2):(1'h1)],
              $signed({reg23, reg94})}));
      for (forvar125 = (1'h0); (forvar125 < (3'h4)); forvar125 = (forvar125 + (1'h1)))
        begin
          reg126 <= (reg102[(3'h6):(2'h2)] ~^ {$unsigned(reg79)});
        end
      reg127 = forvar109[(3'h4):(1'h1)];
    end
  assign wire128 = wire12[(4'h8):(2'h2)];
endmodule
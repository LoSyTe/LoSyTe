(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param931 = ((~&((((7'h43) ? (8'hbd) : (8'hb9)) ^~ (8'hb7)) ? (((8'hb3) || (7'h40)) ? ((7'h40) - (8'h9f)) : (&(7'h43))) : (((8'ha8) | (8'h9f)) >= (+(8'haa))))) >= (((~^(~|(8'hb2))) ? {(+(8'hb1)), (~|(7'h41))} : (((7'h41) | (8'haa)) ? ((8'hba) ? (8'had) : (7'h43)) : {(8'haf)})) ? (((~|(7'h43)) * (&(8'hbd))) < (!{(8'hb5), (8'hb2)})) : (((8'ha4) ? ((8'had) ? (8'ha3) : (7'h40)) : (~(7'h40))) || {{(8'hbc)}, ((8'haa) ^ (8'ha1))}))) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h67b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire0;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire [(4'he):(1'h0)] wire2;
  input wire signed [(4'hc):(1'h0)] wire3;
  input wire [(4'hb):(1'h0)] wire4;
  wire [(5'h13):(1'h0)] wire930;
  wire [(5'h10):(1'h0)] wire929;
  reg signed [(5'h12):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar927 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg926 = (1'h0);
  wire [(5'h12):(1'h0)] wire921;
  reg signed [(3'h5):(1'h0)] reg920 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg919 = (1'h0);
  reg [(4'hd):(1'h0)] reg918 = (1'h0);
  reg [(5'h11):(1'h0)] forvar917 = (1'h0);
  reg [(3'h7):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg915 = (1'h0);
  reg [(3'h4):(1'h0)] reg914 = (1'h0);
  reg [(5'h13):(1'h0)] reg913 = (1'h0);
  reg [(3'h7):(1'h0)] reg912 = (1'h0);
  reg [(5'h10):(1'h0)] forvar911 = (1'h0);
  reg [(4'hb):(1'h0)] reg910 = (1'h0);
  reg [(4'hd):(1'h0)] forvar909 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg908 = (1'h0);
  reg [(5'h13):(1'h0)] reg907 = (1'h0);
  reg [(5'h14):(1'h0)] reg906 = (1'h0);
  reg [(2'h3):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar903 = (1'h0);
  reg [(4'hf):(1'h0)] forvar890 = (1'h0);
  reg [(2'h3):(1'h0)] reg902 = (1'h0);
  reg [(5'h13):(1'h0)] reg901 = (1'h0);
  reg [(4'he):(1'h0)] forvar900 = (1'h0);
  reg [(4'ha):(1'h0)] reg899 = (1'h0);
  reg signed [(4'he):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg897 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg895 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg894 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg893 = (1'h0);
  reg [(2'h3):(1'h0)] reg892 = (1'h0);
  reg [(4'ha):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg890 = (1'h0);
  reg [(4'hf):(1'h0)] reg889 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg888 = (1'h0);
  reg [(4'ha):(1'h0)] reg887 = (1'h0);
  reg [(5'h11):(1'h0)] forvar886 = (1'h0);
  reg [(5'h11):(1'h0)] reg885 = (1'h0);
  reg [(2'h3):(1'h0)] reg884 = (1'h0);
  reg [(5'h11):(1'h0)] reg883 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar882 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg881 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg880 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar879 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg878 = (1'h0);
  reg [(5'h11):(1'h0)] forvar877 = (1'h0);
  wire [(4'he):(1'h0)] wire875;
  reg [(3'h7):(1'h0)] reg5 = (1'h0);
  reg [(5'h14):(1'h0)] reg6 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7 = (1'h0);
  reg [(5'h10):(1'h0)] forvar8 = (1'h0);
  reg [(5'h10):(1'h0)] reg9 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg10 = (1'h0);
  reg [(4'hd):(1'h0)] reg11 = (1'h0);
  reg [(2'h3):(1'h0)] reg12 = (1'h0);
  reg [(4'hc):(1'h0)] reg13 = (1'h0);
  reg [(4'ha):(1'h0)] reg14 = (1'h0);
  reg [(4'hd):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg [(5'h11):(1'h0)] forvar17 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg18 = (1'h0);
  reg [(4'hb):(1'h0)] reg19 = (1'h0);
  reg [(4'h8):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg21 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire816;
  wire signed [(3'h4):(1'h0)] wire818;
  reg signed [(5'h12):(1'h0)] forvar819 = (1'h0);
  reg [(3'h6):(1'h0)] reg820 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg821 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg822 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg823 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg824 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg825 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg819 = (1'h0);
  reg [(5'h11):(1'h0)] forvar820 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar824 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg826 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar827 = (1'h0);
  reg [(2'h2):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg829 = (1'h0);
  reg [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar831 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg832 = (1'h0);
  reg [(5'h12):(1'h0)] reg833 = (1'h0);
  wire [(4'ha):(1'h0)] wire834;
  wire [(3'h4):(1'h0)] wire835;
  reg [(5'h11):(1'h0)] reg836 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire837;
  wire [(4'hc):(1'h0)] wire839;
  reg [(4'hb):(1'h0)] forvar840 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar841 = (1'h0);
  reg [(5'h11):(1'h0)] reg842 = (1'h0);
  reg [(5'h13):(1'h0)] reg843 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg845 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar846 = (1'h0);
  reg [(5'h10):(1'h0)] reg847 = (1'h0);
  reg [(3'h5):(1'h0)] reg848 = (1'h0);
  reg [(4'hb):(1'h0)] reg849 = (1'h0);
  reg [(4'hc):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg851 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar852 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg853 = (1'h0);
  reg [(4'hd):(1'h0)] reg854 = (1'h0);
  reg [(5'h13):(1'h0)] reg855 = (1'h0);
  reg [(5'h10):(1'h0)] reg856 = (1'h0);
  reg [(3'h5):(1'h0)] reg857 = (1'h0);
  reg [(4'hc):(1'h0)] reg858 = (1'h0);
  reg signed [(4'he):(1'h0)] reg859 = (1'h0);
  reg [(5'h15):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar861 = (1'h0);
  reg [(4'hb):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar863 = (1'h0);
  reg [(3'h7):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg867 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar868 = (1'h0);
  reg [(5'h10):(1'h0)] reg869 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg870 = (1'h0);
  reg [(5'h12):(1'h0)] reg871 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg872 = (1'h0);
  wire [(5'h15):(1'h0)] wire873;
  wire [(2'h3):(1'h0)] wire923;
  wire [(5'h15):(1'h0)] wire924;
  assign y = {wire930,
                 wire929,
                 reg928,
                 forvar927,
                 reg926,
                 wire921,
                 reg920,
                 reg919,
                 reg918,
                 forvar917,
                 reg916,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 forvar911,
                 reg910,
                 forvar909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 forvar903,
                 forvar890,
                 reg902,
                 reg901,
                 forvar900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 forvar886,
                 reg885,
                 reg884,
                 reg883,
                 forvar882,
                 reg881,
                 reg880,
                 forvar879,
                 reg878,
                 forvar877,
                 wire875,
                 reg5,
                 reg6,
                 forvar7,
                 forvar8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 forvar17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 wire816,
                 wire818,
                 forvar819,
                 reg820,
                 reg821,
                 reg822,
                 reg823,
                 reg824,
                 reg825,
                 reg819,
                 forvar820,
                 forvar824,
                 reg826,
                 forvar827,
                 reg828,
                 reg829,
                 reg830,
                 forvar831,
                 reg832,
                 reg833,
                 wire834,
                 wire835,
                 reg836,
                 wire837,
                 wire839,
                 forvar840,
                 forvar841,
                 reg842,
                 reg843,
                 reg844,
                 reg845,
                 forvar846,
                 reg847,
                 reg848,
                 reg849,
                 reg850,
                 reg851,
                 forvar852,
                 reg853,
                 reg854,
                 reg855,
                 reg856,
                 reg857,
                 reg858,
                 reg859,
                 reg860,
                 forvar861,
                 reg862,
                 forvar863,
                 reg864,
                 reg865,
                 reg866,
                 reg867,
                 forvar868,
                 reg869,
                 reg870,
                 reg871,
                 reg872,
                 wire873,
                 wire923,
                 wire924,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 = ((wire0 + (wire0 ?
              $unsigned(wire2[(2'h3):(1'h0)]) : $unsigned((!(8'hba))))) ?
          $signed(wire2[(2'h2):(2'h2)]) : wire4[(4'ha):(2'h3)]);
      reg6 = (^$signed(wire2[(2'h2):(1'h1)]));
      for (forvar7 = (1'h0); (forvar7 < (1'h1)); forvar7 = (forvar7 + (1'h1)))
        begin
          for (forvar8 = (1'h0); (forvar8 < (2'h3)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 = (^(reg6[(2'h2):(1'h1)] >= (~|wire4[(3'h5):(3'h5)])));
              reg10 <= wire3;
              reg11 <= reg5;
              reg12 <= wire0[(2'h2):(1'h0)];
            end
          if ((|$unsigned("92Zi68")))
            begin
              reg13 = reg12[(1'h0):(1'h0)];
              reg14 = (|reg6[(3'h5):(1'h1)]);
              reg15 = forvar7;
            end
          else
            begin
              reg13 <= "2uKXT6SiYe";
              reg14 = reg11[(2'h2):(1'h0)];
              reg15 <= (~&$signed((((reg12 ?
                  reg14 : (8'hb0)) ^ (reg12 + wire4)) && (~^$unsigned((8'hb5))))));
              reg16 <= wire4;
            end
          for (forvar17 = (1'h0); (forvar17 < (1'h0)); forvar17 = (forvar17 + (1'h1)))
            begin
              reg18 = $unsigned(wire1[(3'h4):(1'h0)]);
              reg19 = $signed($unsigned((({forvar7} ? wire0 : {reg14, reg10}) ?
                  ((~&reg12) + (reg16 ~^ reg16)) : reg12[(2'h3):(1'h1)])));
              reg20 = $signed($signed($unsigned($unsigned(reg16))));
            end
        end
      reg21 = (8'hb4);
    end
  module22 modinst817 (wire816, clk, wire2, forvar8, reg21, reg13);
  assign wire818 = wire2[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if ((reg10 || {{$unsigned((!wire2)),
              ((forvar17 ^~ (8'hbe)) ? {reg9, wire1} : (wire818 ~^ reg21))}}))
        begin
          for (forvar819 = (1'h0); (forvar819 < (1'h0)); forvar819 = (forvar819 + (1'h1)))
            begin
              reg820 <= $signed(($signed((reg19[(1'h0):(1'h0)] ?
                      forvar7 : ((7'h41) && (8'hb6)))) ?
                  ($signed((forvar8 ? reg21 : reg10)) ?
                      $signed((reg14 ~^ reg19)) : $signed(reg19[(1'h1):(1'h0)])) : $unsigned(((^~(8'haa)) * reg19[(4'ha):(4'ha)]))));
              reg821 = $unsigned(reg820);
              reg822 = forvar17[(4'h8):(1'h1)];
              reg823 <= ($unsigned(("6YTaLvpze" < (wire0[(2'h3):(2'h3)] ?
                      reg9 : (reg20 <= forvar8)))) ?
                  ((|($signed(wire2) ? $unsigned((8'ha4)) : (|(8'hb9)))) ?
                      $signed(reg9) : reg821[(1'h1):(1'h1)]) : $signed((^~$signed(((8'h9c) << forvar8)))));
            end
          if ((-(reg19 ^~ $unsigned($unsigned($signed(reg6))))))
            begin
              reg824 = $unsigned(((((reg9 < wire818) ?
                      (forvar819 ? wire4 : forvar17) : (reg16 ?
                          (8'ha2) : (8'hbf))) <<< ($unsigned((7'h41)) ?
                      $signed(reg14) : $signed(reg12))) ?
                  $unsigned({$signed(reg16)}) : $signed($signed(reg18))));
              reg825 = {wire1};
            end
          else
            begin
              reg824 = (({reg19[(2'h2):(2'h2)], $signed("")} ?
                  (^~{$unsigned(reg16),
                      "EQXtQ4Pio6LJVidU"}) : reg16[(3'h6):(2'h3)]) >= ($signed(({reg15} ^ $signed(reg16))) ?
                  {$signed((reg13 ?
                          reg12 : reg13))} : (forvar17[(1'h0):(1'h0)] >= $signed("J"))));
            end
        end
      else
        begin
          reg819 <= $unsigned({(!forvar8[(4'hd):(3'h6)])});
          for (forvar820 = (1'h0); (forvar820 < (2'h3)); forvar820 = (forvar820 + (1'h1)))
            begin
              reg821 <= $unsigned(reg13[(2'h2):(1'h0)]);
              reg822 <= {$unsigned(reg6[(5'h12):(5'h10)])};
            end
          reg823 <= $unsigned(reg5);
          for (forvar824 = (1'h0); (forvar824 < (3'h4)); forvar824 = (forvar824 + (1'h1)))
            begin
              reg825 = (($signed($signed((|reg823))) ^~ (!$signed((wire1 ?
                  reg16 : reg14)))) > ((!($signed(wire818) ?
                  (reg5 ?
                      reg819 : reg16) : (~^reg825))) ~^ ($signed(reg823[(3'h5):(3'h4)]) ~^ reg18[(2'h2):(2'h2)])));
            end
        end
      reg826 <= ((-reg820) <<< forvar820);
      for (forvar827 = (1'h0); (forvar827 < (2'h2)); forvar827 = (forvar827 + (1'h1)))
        begin
          if ({((-{{forvar17, reg824}}) ^~ (forvar820 ?
                  (!$unsigned(reg11)) : ((reg11 >> wire4) & (~|(8'h9d)))))})
            begin
              reg828 = $signed(((!(+$unsigned(reg6))) && (|$signed($unsigned(wire4)))));
              reg829 <= ({$signed(((8'ha5) ? (reg824 == (8'hb6)) : reg824)),
                  ((forvar8[(4'h9):(4'h9)] ?
                      (reg20 ?
                          (8'hbc) : (8'ha9)) : {reg820}) << (wire3[(1'h0):(1'h0)] && $signed(reg824)))} != reg823);
              reg830 <= ($signed((~|$signed({wire3}))) ?
                  $unsigned((reg819[(2'h2):(1'h1)] ?
                      {reg825,
                          $unsigned((8'hbb))} : reg6[(4'hd):(4'hd)])) : (reg21 ?
                      reg19[(3'h6):(3'h6)] : (((|reg828) ?
                              {reg819} : (forvar824 ? reg18 : reg6)) ?
                          $signed((reg828 ?
                              wire3 : reg16)) : ((&forvar827) || (reg11 << forvar820)))));
            end
          else
            begin
              reg828 = $unsigned(reg820[(1'h0):(1'h0)]);
              reg829 <= forvar819;
            end
          for (forvar831 = (1'h0); (forvar831 < (2'h2)); forvar831 = (forvar831 + (1'h1)))
            begin
              reg832 <= $unsigned(($signed(((reg12 == (8'hab)) + {(7'h40)})) >= reg10[(3'h6):(3'h5)]));
            end
        end
      reg833 = (~$signed($unsigned(reg6[(4'ha):(2'h2)])));
    end
  assign wire834 = $unsigned(wire2);
  assign wire835 = reg20;
  always
    @(posedge clk) begin
      reg836 = (~^reg829[(5'h10):(5'h10)]);
    end
  module204 modinst838 (.wire207(wire816), .wire206(forvar819), .wire205(forvar824), .clk(clk), .y(wire837), .wire208(reg829));
  assign wire839 = forvar831[(4'h9):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar840 = (1'h0); (forvar840 < (3'h4)); forvar840 = (forvar840 + (1'h1)))
        begin
          for (forvar841 = (1'h0); (forvar841 < (2'h3)); forvar841 = (forvar841 + (1'h1)))
            begin
              reg842 = reg6;
              reg843 <= ($signed({reg822,
                  forvar819[(2'h3):(2'h3)]}) ^~ ((($signed(reg19) && (&forvar841)) > $signed($unsigned(reg823))) ?
                  (($signed(wire818) ? (|reg15) : reg18[(3'h6):(1'h1)]) ?
                      $unsigned("wHxS") : $unsigned((reg19 ?
                          (8'hba) : reg5))) : (reg6[(3'h4):(3'h4)] ?
                      (((8'hba) == forvar831) ?
                          forvar819 : wire818) : $signed((reg832 ?
                          forvar841 : wire839)))));
              reg844 <= ("vHwWrfqeOzwt" ?
                  {(~(+$unsigned(reg820))),
                      $unsigned((reg828[(1'h0):(1'h0)] ?
                          (&reg14) : $signed(reg16)))} : (8'hac));
              reg845 <= (wire3[(4'ha):(4'ha)] >> $unsigned(forvar819[(3'h7):(3'h6)]));
            end
          for (forvar846 = (1'h0); (forvar846 < (1'h1)); forvar846 = (forvar846 + (1'h1)))
            begin
              reg847 <= wire0[(4'h8):(1'h1)];
              reg848 = ("YL66IvnzMmR0LSN" ?
                  ({((8'hbb) ?
                          {reg10} : reg819[(1'h0):(1'h0)])} ^~ reg830) : reg843[(3'h7):(3'h6)]);
              reg849 = reg16[(1'h1):(1'h1)];
              reg850 = (~&(^reg21[(5'h12):(2'h2)]));
              reg851 <= (~^$unsigned(($signed(reg14[(2'h2):(1'h1)]) ?
                  $unsigned({(8'h9d), reg20}) : forvar17[(3'h5):(1'h1)])));
            end
          for (forvar852 = (1'h0); (forvar852 < (1'h1)); forvar852 = (forvar852 + (1'h1)))
            begin
              reg853 = {$signed(($signed((forvar841 & reg14)) ?
                      (reg6[(4'hd):(4'h8)] ? (~|forvar831) : reg833) : reg822)),
                  ((|(8'ha5)) < reg20[(1'h0):(1'h0)])};
            end
          if ($signed((!(wire839[(1'h1):(1'h0)] ?
              ($unsigned(reg5) ^ wire837[(3'h5):(2'h3)]) : ($unsigned(reg836) << (forvar831 ?
                  reg12 : reg6))))))
            begin
              reg854 <= ($unsigned({forvar831}) ?
                  {(~|($unsigned(reg845) ~^ {reg825, reg828})),
                      reg853} : wire835[(2'h2):(1'h0)]);
            end
          else
            begin
              reg854 <= reg853[(3'h4):(1'h0)];
              reg855 <= (($unsigned((~&forvar852[(1'h0):(1'h0)])) ?
                  $unsigned(((forvar824 != wire3) != (~|forvar820))) : reg849[(4'hb):(4'h9)]) && ($unsigned($unsigned((forvar7 ?
                  reg832 : wire834))) >= reg11));
              reg856 = reg20;
              reg857 <= $unsigned(({(forvar17 <<< (+reg16)), $signed(reg855)} ?
                  (~reg829) : $unsigned("kY1Skkk")));
            end
          reg858 = ((reg830 ?
              $signed($unsigned((forvar819 >= reg828))) : $signed($signed((reg825 ?
                  reg5 : (8'ha4))))) & (~&""));
        end
      reg859 = (reg16 * reg853[(2'h3):(2'h2)]);
      reg860 = wire835;
      for (forvar861 = (1'h0); (forvar861 < (2'h3)); forvar861 = (forvar861 + (1'h1)))
        begin
          reg862 = (8'hb0);
          for (forvar863 = (1'h0); (forvar863 < (1'h1)); forvar863 = (forvar863 + (1'h1)))
            begin
              reg864 = "q0fFZ9i7nYZ";
              reg865 = (($signed($unsigned("84nS")) ?
                  $signed(({forvar17,
                      reg9} <<< (wire3 & reg829))) : $unsigned($signed(((8'hb7) ~^ reg844)))) <<< (-reg858));
              reg866 <= ($signed((((-wire816) ?
                      $signed(reg823) : $signed(forvar852)) >= ({wire837} ?
                      $signed(reg10) : (8'ha6)))) ?
                  $signed($signed(((reg842 + reg821) > (reg6 ~^ reg862)))) : reg823[(3'h5):(2'h3)]);
            end
          reg867 = $signed({$signed((+forvar846[(2'h3):(2'h3)]))});
          for (forvar868 = (1'h0); (forvar868 < (2'h3)); forvar868 = (forvar868 + (1'h1)))
            begin
              reg869 <= "7VbfZ1";
              reg870 <= reg829;
              reg871 = reg18;
              reg872 <= ((8'hb4) ?
                  forvar7 : $signed($unsigned($unsigned({wire2, reg842}))));
            end
        end
    end
  module326 modinst874 (wire873, clk, reg872, reg848, forvar8, reg20, reg860);
  module204 modinst876 (wire875, clk, forvar17, reg844, forvar841, reg819);
  always
    @(posedge clk) begin
      for (forvar877 = (1'h0); (forvar877 < (3'h4)); forvar877 = (forvar877 + (1'h1)))
        begin
          reg878 <= forvar841;
        end
      for (forvar879 = (1'h0); (forvar879 < (3'h4)); forvar879 = (forvar879 + (1'h1)))
        begin
          if (((reg856[(1'h1):(1'h1)] ^ reg6[(4'he):(2'h2)]) - (-((-{(8'hae),
              reg829}) & $signed(wire2)))))
            begin
              reg880 = (8'haa);
            end
          else
            begin
              reg880 = ((reg822[(2'h3):(2'h2)] ?
                  $unsigned($unsigned((^~wire873))) : wire834[(4'ha):(3'h5)]) || wire837[(4'h8):(1'h0)]);
              reg881 <= (reg864 ? forvar868 : $unsigned(reg16));
            end
          for (forvar882 = (1'h0); (forvar882 < (1'h1)); forvar882 = (forvar882 + (1'h1)))
            begin
              reg883 = $unsigned($unsigned($signed(forvar7[(4'hd):(4'ha)])));
              reg884 <= $unsigned($unsigned(wire2[(4'ha):(3'h4)]));
              reg885 <= reg21;
            end
          for (forvar886 = (1'h0); (forvar886 < (1'h0)); forvar886 = (forvar886 + (1'h1)))
            begin
              reg887 = $signed($signed($signed((wire1[(1'h0):(1'h0)] ?
                  (reg843 == wire835) : reg819))));
              reg888 <= $unsigned((^~"WvxqPRq"));
            end
          reg889 <= ($unsigned(reg888) ? (~&{reg880[(3'h7):(3'h4)]}) : reg885);
        end
      if ($unsigned((|((~&(reg855 ~^ reg12)) > {(&reg853)}))))
        begin
          if (((wire2 << ((^~"FwrcQSxDUT98") != ({reg888} != {reg822}))) | forvar882))
            begin
              reg890 = $signed($signed(reg864));
              reg891 = $signed(((reg872 ?
                      (reg884 ? {reg836} : "gpHPn1") : (|(!reg11))) ?
                  ({((8'hae) ? reg845 : reg842), $unsigned(reg10)} ?
                      $signed($signed(forvar846)) : (8'ha0)) : (reg824[(3'h4):(1'h1)] ?
                      $unsigned(reg888) : reg883[(4'hb):(4'h8)])));
              reg892 <= forvar819;
              reg893 = (&forvar868[(2'h3):(2'h2)]);
            end
          else
            begin
              reg890 <= $unsigned($signed(($unsigned(reg860[(5'h10):(1'h1)]) ?
                  reg866[(4'he):(2'h2)] : $unsigned((~&reg19)))));
              reg891 <= reg14;
              reg892 = $signed((reg12[(1'h1):(1'h1)] ^~ (($signed(reg884) == reg823) ?
                  ((reg11 ? reg891 : (8'hb9)) << $signed((8'h9f))) : {(wire837 ?
                          forvar17 : forvar819),
                      {reg869}})));
              reg893 = (((forvar17[(3'h5):(2'h3)] || (~^((8'hb0) ?
                      reg845 : forvar863))) && $signed(wire816)) ?
                  {((|$unsigned(forvar852)) ~^ (|$unsigned(reg880)))} : $unsigned(reg847[(4'h9):(3'h5)]));
            end
          if ((reg885 ?
              (reg824[(1'h1):(1'h1)] ?
                  ({reg880} > $signed((~reg892))) : (^$unsigned((!(8'ha7))))) : $signed($unsigned(({reg854} ?
                  $unsigned((8'ha4)) : $signed(reg850))))))
            begin
              reg894 <= wire4;
              reg895 = $signed($signed(((8'haa) || (~|(8'h9d)))));
              reg896 = (|forvar8[(4'hb):(3'h4)]);
              reg897 = $signed($signed($signed($unsigned($unsigned(reg829)))));
              reg898 <= reg819[(3'h7):(1'h0)];
            end
          else
            begin
              reg894 <= $signed("WVm94ETkfAxKMZOXyONw");
              reg895 = $signed($signed((&{(forvar841 & reg885),
                  wire837[(4'ha):(1'h0)]})));
              reg896 = (&("9BxzionAyE1xCE43mmR" <<< reg832));
              reg897 <= "Tw4g4Wq";
            end
          reg899 <= $signed(((^~(reg869[(4'hd):(3'h7)] | {(8'hb2)})) ?
              {{$unsigned(reg15), $unsigned(reg884)}} : reg858));
          for (forvar900 = (1'h0); (forvar900 < (2'h3)); forvar900 = (forvar900 + (1'h1)))
            begin
              reg901 = $signed($unsigned(($unsigned($signed(wire4)) < (~|forvar7))));
              reg902 = (reg843[(5'h11):(4'hc)] ? reg869 : wire1);
            end
        end
      else
        begin
          for (forvar890 = (1'h0); (forvar890 < (3'h4)); forvar890 = (forvar890 + (1'h1)))
            begin
              reg891 <= ((wire3[(4'hc):(3'h5)] ?
                      (|$signed($unsigned(reg844))) : (&(!(forvar17 ?
                          reg819 : (8'haf))))) ?
                  reg853[(1'h0):(1'h0)] : (8'hb6));
            end
          reg892 = (&{(^$unsigned($unsigned(forvar8)))});
        end
      for (forvar903 = (1'h0); (forvar903 < (3'h4)); forvar903 = (forvar903 + (1'h1)))
        begin
          reg904 <= $signed({$signed(((reg822 || (8'had)) <= reg19[(2'h2):(1'h1)]))});
          if (($signed($unsigned((~$unsigned(reg5)))) - (forvar824[(2'h3):(1'h0)] == forvar882[(2'h3):(1'h1)])))
            begin
              reg905 <= {$signed(reg883[(3'h6):(2'h3)]),
                  ($signed({(reg894 ^ reg895),
                      (~&(8'ha8))}) && (($unsigned(reg842) ?
                      reg899[(3'h4):(1'h1)] : wire834[(2'h2):(1'h0)]) & $unsigned(forvar820)))};
              reg906 <= $signed($signed($unsigned((8'h9c))));
              reg907 = reg862[(3'h7):(2'h2)];
              reg908 = $unsigned({{reg11}});
            end
          else
            begin
              reg905 = $signed("sC");
              reg906 <= $signed(forvar861);
            end
          for (forvar909 = (1'h0); (forvar909 < (2'h3)); forvar909 = (forvar909 + (1'h1)))
            begin
              reg910 <= wire2;
            end
          for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
            begin
              reg912 = "sPwuXOioPN8wIKxq";
              reg913 <= ($signed(({(reg869 ? reg21 : reg14),
                      $unsigned(reg850)} ?
                  forvar909 : ((reg894 ?
                      forvar886 : reg895) >= reg10))) << $signed($signed((~|reg10[(1'h0):(1'h0)]))));
              reg914 <= reg894;
              reg915 <= (8'ha0);
              reg916 = ($signed(((~|(8'hab)) ?
                      reg9 : $signed((reg845 - reg898)))) ?
                  ((~&($unsigned(reg865) || (reg862 ?
                      (7'h40) : reg878))) ^~ (&{(^~(8'hbf))})) : forvar900[(4'hc):(3'h6)]);
            end
          for (forvar917 = (1'h0); (forvar917 < (2'h2)); forvar917 = (forvar917 + (1'h1)))
            begin
              reg918 <= $signed((&(~reg823)));
              reg919 <= reg899;
              reg920 = $unsigned((reg844 * (!$unsigned((wire1 ?
                  (8'hbc) : reg878)))));
            end
        end
    end
  module27 modinst922 (wire921, clk, forvar877, reg883, wire875, reg830, forvar886);
  assign wire923 = (reg880[(2'h3):(1'h0)] ?
                       $signed((~&reg897[(4'ha):(4'ha)])) : {(~|(8'ha1)),
                           {$signed((^~forvar868)), wire2}});
  module326 modinst925 (.wire328(reg825), .clk(clk), .wire327(wire837), .wire330(reg910), .y(wire924), .wire331(reg907), .wire329(reg894));
  always
    @(posedge clk) begin
      reg926 <= $unsigned(($unsigned($unsigned(forvar819[(4'hc):(3'h4)])) ?
          reg856 : {$unsigned(reg880), ($unsigned(reg844) * (~^reg828))}));
      for (forvar927 = (1'h0); (forvar927 < (1'h0)); forvar927 = (forvar927 + (1'h1)))
        begin
          reg928 <= {$unsigned(forvar17), $signed(wire835[(1'h0):(1'h0)])};
        end
    end
  assign wire929 = {(reg905 ?
                           ("EZz6gZE" ?
                               (~|(~&reg896)) : forvar819[(5'h10):(3'h4)]) : $unsigned(forvar819[(4'h8):(1'h0)]))};
  assign wire930 = reg855[(5'h13):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module22  (y, clk, wire26, wire25, wire24, wire23);
  output wire [(32'h888):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire26;
  input wire [(4'he):(1'h0)] wire25;
  input wire [(5'h14):(1'h0)] wire24;
  input wire [(4'h8):(1'h0)] wire23;
  reg [(4'h9):(1'h0)] reg812 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg815 = (1'h0);
  reg [(2'h3):(1'h0)] reg814 = (1'h0);
  reg [(4'hb):(1'h0)] reg813 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar812 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg811 = (1'h0);
  reg [(4'hd):(1'h0)] reg810 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar809 = (1'h0);
  reg [(5'h12):(1'h0)] forvar791 = (1'h0);
  reg [(4'ha):(1'h0)] reg808 = (1'h0);
  reg [(5'h15):(1'h0)] reg807 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg806 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg805 = (1'h0);
  reg [(4'hf):(1'h0)] reg804 = (1'h0);
  reg [(5'h11):(1'h0)] reg803 = (1'h0);
  reg signed [(4'he):(1'h0)] reg802 = (1'h0);
  reg [(4'h8):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg799 = (1'h0);
  reg [(5'h15):(1'h0)] reg798 = (1'h0);
  reg [(4'h9):(1'h0)] reg797 = (1'h0);
  reg [(4'he):(1'h0)] forvar796 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg795 = (1'h0);
  reg [(5'h12):(1'h0)] reg794 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg793 = (1'h0);
  reg [(4'hf):(1'h0)] reg792 = (1'h0);
  reg signed [(4'he):(1'h0)] reg791 = (1'h0);
  reg [(5'h11):(1'h0)] reg790 = (1'h0);
  reg [(4'h9):(1'h0)] reg789 = (1'h0);
  reg [(3'h7):(1'h0)] reg788 = (1'h0);
  reg [(3'h6):(1'h0)] reg787 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar786 = (1'h0);
  reg [(4'h9):(1'h0)] reg785 = (1'h0);
  reg signed [(4'he):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg783 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg782 = (1'h0);
  reg [(4'hd):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg780 = (1'h0);
  reg [(3'h5):(1'h0)] reg779 = (1'h0);
  reg [(5'h12):(1'h0)] reg778 = (1'h0);
  reg [(3'h5):(1'h0)] forvar777 = (1'h0);
  reg [(3'h6):(1'h0)] reg776 = (1'h0);
  reg [(5'h12):(1'h0)] forvar775 = (1'h0);
  reg [(4'ha):(1'h0)] reg774 = (1'h0);
  reg [(4'h8):(1'h0)] reg773 = (1'h0);
  reg [(5'h15):(1'h0)] reg772 = (1'h0);
  reg [(4'hd):(1'h0)] reg771 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg770 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar769 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg767 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar766 = (1'h0);
  reg [(4'h8):(1'h0)] reg765 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg764 = (1'h0);
  reg [(5'h10):(1'h0)] forvar763 = (1'h0);
  reg [(3'h4):(1'h0)] forvar762 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg760 = (1'h0);
  wire [(4'hb):(1'h0)] wire755;
  wire [(3'h5):(1'h0)] wire754;
  wire signed [(5'h10):(1'h0)] wire753;
  wire signed [(4'hc):(1'h0)] wire752;
  reg [(2'h3):(1'h0)] reg751 = (1'h0);
  reg [(4'he):(1'h0)] reg750 = (1'h0);
  reg [(5'h15):(1'h0)] reg749 = (1'h0);
  reg [(4'hd):(1'h0)] reg748 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg747 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg746 = (1'h0);
  reg [(5'h14):(1'h0)] reg745 = (1'h0);
  reg [(2'h2):(1'h0)] forvar744 = (1'h0);
  reg [(5'h11):(1'h0)] forvar743 = (1'h0);
  reg [(4'hd):(1'h0)] reg742 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg741 = (1'h0);
  reg [(5'h15):(1'h0)] reg740 = (1'h0);
  reg [(3'h5):(1'h0)] reg739 = (1'h0);
  reg [(3'h7):(1'h0)] forvar738 = (1'h0);
  reg [(2'h3):(1'h0)] reg737 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg736 = (1'h0);
  reg [(4'ha):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg734 = (1'h0);
  reg [(5'h10):(1'h0)] reg733 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar732 = (1'h0);
  reg [(3'h7):(1'h0)] reg731 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg729 = (1'h0);
  reg [(5'h12):(1'h0)] reg728 = (1'h0);
  reg [(4'ha):(1'h0)] reg727 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar726 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg725 = (1'h0);
  reg [(5'h14):(1'h0)] reg724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg723 = (1'h0);
  reg [(3'h5):(1'h0)] reg722 = (1'h0);
  reg [(5'h12):(1'h0)] forvar721 = (1'h0);
  reg [(5'h11):(1'h0)] reg720 = (1'h0);
  reg [(3'h7):(1'h0)] reg719 = (1'h0);
  reg [(5'h14):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg716 = (1'h0);
  reg [(5'h12):(1'h0)] reg715 = (1'h0);
  reg [(4'h8):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg713 = (1'h0);
  reg [(5'h15):(1'h0)] reg712 = (1'h0);
  reg [(5'h11):(1'h0)] forvar711 = (1'h0);
  reg [(5'h12):(1'h0)] reg711 = (1'h0);
  reg [(4'h8):(1'h0)] reg710 = (1'h0);
  reg [(5'h14):(1'h0)] reg709 = (1'h0);
  reg [(5'h15):(1'h0)] reg708 = (1'h0);
  reg [(4'ha):(1'h0)] reg707 = (1'h0);
  reg [(2'h2):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar705 = (1'h0);
  reg [(3'h7):(1'h0)] reg704 = (1'h0);
  reg [(4'ha):(1'h0)] forvar703 = (1'h0);
  reg [(3'h5):(1'h0)] reg702 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg701 = (1'h0);
  reg [(5'h13):(1'h0)] reg700 = (1'h0);
  reg [(2'h2):(1'h0)] reg699 = (1'h0);
  reg [(3'h6):(1'h0)] forvar698 = (1'h0);
  reg [(2'h3):(1'h0)] reg697 = (1'h0);
  reg [(4'ha):(1'h0)] forvar696 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg695 = (1'h0);
  reg [(4'hf):(1'h0)] forvar694 = (1'h0);
  reg [(3'h5):(1'h0)] reg693 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire692;
  reg signed [(2'h3):(1'h0)] reg691 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg690 = (1'h0);
  reg [(4'hc):(1'h0)] reg689 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg688 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg687 = (1'h0);
  reg [(3'h4):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg685 = (1'h0);
  reg [(5'h12):(1'h0)] forvar684 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg683 = (1'h0);
  reg [(4'h8):(1'h0)] forvar679 = (1'h0);
  reg [(4'h8):(1'h0)] reg682 = (1'h0);
  reg [(5'h14):(1'h0)] reg681 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg680 = (1'h0);
  reg [(3'h6):(1'h0)] reg679 = (1'h0);
  reg [(5'h12):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar677 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire383;
  wire [(4'he):(1'h0)] wire325;
  wire signed [(5'h15):(1'h0)] wire324;
  wire signed [(5'h11):(1'h0)] wire323;
  wire [(4'h8):(1'h0)] wire322;
  wire signed [(4'hc):(1'h0)] wire320;
  reg [(3'h4):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg203 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg202 = (1'h0);
  reg [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(5'h11):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar199 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar195 = (1'h0);
  reg [(4'hb):(1'h0)] forvar192 = (1'h0);
  reg [(4'hb):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  reg [(2'h2):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg191 = (1'h0);
  reg [(4'hb):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg189 = (1'h0);
  reg [(5'h14):(1'h0)] forvar188 = (1'h0);
  reg [(4'he):(1'h0)] forvar187 = (1'h0);
  reg [(4'h9):(1'h0)] reg186 = (1'h0);
  reg [(3'h7):(1'h0)] reg185 = (1'h0);
  reg [(5'h15):(1'h0)] reg184 = (1'h0);
  reg [(4'hc):(1'h0)] reg183 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg [(3'h5):(1'h0)] forvar181 = (1'h0);
  reg [(2'h2):(1'h0)] forvar180 = (1'h0);
  reg [(4'he):(1'h0)] reg179 = (1'h0);
  reg [(4'hf):(1'h0)] reg178 = (1'h0);
  reg [(5'h13):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg176 = (1'h0);
  reg [(5'h10):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg174 = (1'h0);
  reg [(3'h6):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] forvar171 = (1'h0);
  wire [(5'h10):(1'h0)] wire169;
  wire [(4'hd):(1'h0)] wire675;
  wire [(3'h6):(1'h0)] wire757;
  wire [(5'h11):(1'h0)] wire758;
  assign y = {reg812,
                 reg815,
                 reg814,
                 reg813,
                 forvar812,
                 reg811,
                 reg810,
                 forvar809,
                 forvar791,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 forvar796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg787,
                 forvar786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 forvar777,
                 reg776,
                 forvar775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 forvar769,
                 reg768,
                 reg767,
                 forvar766,
                 reg765,
                 reg764,
                 forvar763,
                 forvar762,
                 reg761,
                 reg760,
                 wire755,
                 wire754,
                 wire753,
                 wire752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 forvar744,
                 forvar743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 forvar738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 forvar732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 forvar726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 forvar721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 forvar711,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 forvar705,
                 reg704,
                 forvar703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 forvar698,
                 reg697,
                 forvar696,
                 reg695,
                 forvar694,
                 reg693,
                 wire692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 forvar684,
                 reg683,
                 forvar679,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 forvar677,
                 wire383,
                 wire325,
                 wire324,
                 wire323,
                 wire322,
                 wire320,
                 reg199,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 forvar199,
                 forvar195,
                 forvar192,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 forvar188,
                 forvar187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 forvar181,
                 forvar180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 forvar171,
                 wire169,
                 wire675,
                 wire757,
                 wire758,
                 (1'h0)};
  module27 modinst170 (.wire31(wire25), .clk(clk), .wire28((8'haa)), .wire32(wire23), .wire30(wire26), .y(wire169), .wire29(wire24));
  always
    @(posedge clk) begin
      for (forvar171 = (1'h0); (forvar171 < (2'h3)); forvar171 = (forvar171 + (1'h1)))
        begin
          reg172 <= $signed(($signed(wire169) ?
              ((wire25[(1'h1):(1'h0)] << wire26[(4'h8):(3'h5)]) == (wire24 ?
                  (wire23 ?
                      (8'ha1) : forvar171) : $signed(wire25))) : $unsigned("dB6MmEoNHBO9of9NzN")));
          reg173 = (8'hbe);
          reg174 <= $unsigned(((((reg173 <<< reg173) ?
                  {(8'ha7), wire24} : reg173) + wire169[(2'h2):(1'h0)]) ?
              (~"DD") : ($signed(reg173) ?
                  (forvar171 <<< ((8'hb1) <= reg173)) : ((reg173 ?
                      forvar171 : reg172) == reg173[(3'h4):(2'h2)]))));
          if (($signed(((!forvar171) >> wire24)) ?
              (+wire169) : (-$unsigned(({(8'hb6), forvar171} ?
                  (8'hb6) : {(8'ha3)})))))
            begin
              reg175 = (7'h40);
              reg176 <= ({reg173[(2'h2):(2'h2)]} ~^ (|((|$unsigned(reg172)) ?
                  forvar171[(5'h15):(5'h12)] : (((8'hb0) & reg173) ?
                      {wire25, reg175} : ((8'hae) ? wire25 : (8'hbe))))));
              reg177 <= {wire23, $unsigned(((8'h9d) < reg172[(3'h5):(3'h5)]))};
              reg178 <= {{$signed(($unsigned(reg172) + reg172)), reg174},
                  $unsigned(wire23[(4'h8):(2'h3)])};
              reg179 = $signed((!(8'hb6)));
            end
          else
            begin
              reg175 = wire24;
              reg176 <= (wire169[(3'h7):(2'h3)] ?
                  reg174 : $unsigned((!$signed(wire24))));
              reg177 <= reg175[(4'hd):(4'hc)];
              reg178 = $signed("wOdcNeMviZORRVqwlaqN");
            end
        end
      for (forvar180 = (1'h0); (forvar180 < (2'h2)); forvar180 = (forvar180 + (1'h1)))
        begin
          for (forvar181 = (1'h0); (forvar181 < (3'h4)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 = (wire23 ?
                  $unsigned(forvar171) : {(^~forvar181), (8'haa)});
              reg183 <= (&("zQhOZp" || $unsigned((&wire23[(3'h7):(1'h1)]))));
              reg184 = (~{$unsigned(wire25),
                  $unsigned({reg174[(2'h3):(1'h0)]})});
              reg185 <= {($unsigned($signed(reg182)) ?
                      (({reg172} | wire23) ?
                          wire169[(4'hf):(4'hf)] : $unsigned($signed(wire26))) : ($signed(wire23[(4'h8):(4'h8)]) ?
                          $signed($signed(reg174)) : $signed((reg175 ?
                              reg174 : reg174)))),
                  $unsigned((wire25[(1'h1):(1'h0)] ?
                      (reg179 ? wire169 : $signed(reg184)) : $unsigned({reg177,
                          wire25})))};
              reg186 <= ((~^$signed(((reg183 >>> reg179) ?
                      (|wire24) : wire26))) ?
                  (((~&$signed(reg185)) ^ reg185) ?
                      $signed(reg178[(2'h3):(1'h0)]) : (!(8'ha1))) : $unsigned($unsigned(wire26)));
            end
        end
      for (forvar187 = (1'h0); (forvar187 < (1'h1)); forvar187 = (forvar187 + (1'h1)))
        begin
          for (forvar188 = (1'h0); (forvar188 < (3'h4)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= (~^forvar188);
              reg190 <= {((~reg186[(3'h6):(3'h4)]) ?
                      $unsigned($signed($signed(forvar187))) : (reg182 ?
                          reg173 : ($unsigned((8'hb8)) - $signed(reg184)))),
                  (reg177[(2'h3):(1'h0)] ?
                      reg185[(3'h6):(1'h1)] : (&reg182[(2'h2):(2'h2)]))};
            end
          reg191 <= wire169;
        end
      if (wire26)
        begin
          if ($signed((reg189[(5'h12):(5'h10)] ?
              wire25[(4'h9):(1'h0)] : reg191)))
            begin
              reg192 = $signed(reg183[(4'h9):(3'h6)]);
              reg193 <= (&forvar187[(2'h2):(1'h0)]);
              reg194 = {(reg176 >= $signed((^$signed(reg190)))),
                  $unsigned($unsigned($unsigned($signed((8'hbf)))))};
            end
          else
            begin
              reg192 <= {$unsigned((~&(~^(~&reg178)))),
                  {$signed((forvar187 ?
                          (forvar180 ? reg182 : wire25) : (!reg182))),
                      (&(((8'ha1) * reg179) ? (^~(8'hb6)) : (^~forvar171)))}};
              reg193 <= (~&((forvar187[(2'h2):(2'h2)] ?
                  ($unsigned(wire25) ?
                      ((8'hb1) ?
                          forvar180 : reg184) : reg189) : reg194[(3'h4):(3'h4)]) != ($unsigned($signed(forvar180)) & $signed((~&forvar188)))));
              reg194 <= (|$signed(($signed(reg175) >> reg183)));
              reg195 <= reg178;
              reg196 = "ksysv";
            end
          reg197 = (8'ha7);
          reg198 = reg174;
        end
      else
        begin
          for (forvar192 = (1'h0); (forvar192 < (2'h3)); forvar192 = (forvar192 + (1'h1)))
            begin
              reg193 <= (((reg196 ?
                      reg176[(1'h1):(1'h1)] : $signed(forvar188)) > (8'h9e)) ?
                  (~((|((8'hb2) ^~ reg189)) <<< $unsigned((+reg194)))) : reg196[(4'hb):(3'h4)]);
              reg194 = $unsigned(((((!forvar180) << $unsigned(forvar188)) ?
                  {(reg197 ?
                          wire25 : (8'hb5))} : {$unsigned(reg191)}) < ($unsigned(reg192[(2'h3):(1'h1)]) ?
                  ($unsigned(reg197) ^ $unsigned(wire24)) : ((reg179 >> forvar181) ?
                      (~|reg198) : reg191[(5'h10):(4'ha)]))));
            end
          for (forvar195 = (1'h0); (forvar195 < (2'h2)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 <= ((forvar192[(3'h7):(3'h4)] ?
                  (-((reg186 ?
                      forvar180 : forvar181) & reg182)) : reg179) ^~ (8'hbe));
              reg197 = "ynw8f2LuM";
            end
          reg198 = ((($unsigned((~^forvar187)) ?
                  (forvar195 >>> ((8'hb1) ^ reg192)) : {(!reg195)}) ?
              ($signed({wire169, (8'had)}) ?
                  (&(~|reg189)) : ((8'hb0) ?
                      $unsigned(reg196) : (wire169 ?
                          reg196 : reg177))) : $signed((~|(&reg193)))) != reg184);
        end
    end
  always
    @(posedge clk) begin
      if (($unsigned($unsigned(($signed(reg194) < $unsigned(forvar187)))) ?
          $signed(((8'ha7) & (^(reg195 ^ forvar195)))) : reg192))
        begin
          for (forvar199 = (1'h0); (forvar199 < (2'h3)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 = ($unsigned({reg194[(3'h5):(3'h4)], (|(|reg173))}) ?
                  (($signed(reg197) == (!$signed((8'had)))) & (reg178 ?
                      (!((8'ha9) >> reg189)) : (&$signed(forvar192)))) : forvar171);
              reg201 = reg184;
              reg202 <= (!$unsigned($unsigned($unsigned((^reg179)))));
              reg203 = (~$unsigned(reg191[(4'h9):(4'h8)]));
            end
        end
      else
        begin
          reg199 = {(^~"IN8"),
              (reg189[(4'h9):(3'h5)] ?
                  ($signed(wire25) ^~ (&$signed(wire169))) : ({$unsigned(reg183)} != (8'hb3)))};
        end
    end
  module204 modinst321 (.wire205(wire24), .clk(clk), .y(wire320), .wire206(forvar188), .wire207(reg200), .wire208(reg196));
  assign wire322 = $signed((($signed($unsigned(reg176)) ^~ "kKf0JLRGvLdO6u091c") ?
                       $signed($signed((reg193 << wire26))) : $signed(forvar195)));
  assign wire323 = $signed((reg203[(3'h6):(1'h1)] ?
                       ("POz35n1AZM0" ?
                           (~^(^forvar199)) : {(reg185 ?
                                   reg193 : wire322)}) : (forvar171[(5'h11):(2'h2)] ?
                           $signed($unsigned(reg174)) : (|$unsigned(reg186)))));
  assign wire324 = reg202;
  assign wire325 = ($signed(("HpJP3ZzlAfulUvulm7YD" > $signed(reg198[(4'h8):(1'h1)]))) ?
                       (8'haa) : wire25);
  module326 modinst384 (wire383, clk, forvar171, wire323, wire169, wire26, forvar181);
  module385 modinst676 (.wire386(reg190), .wire389(reg203), .wire387(wire25), .wire390(forvar171), .y(wire675), .clk(clk), .wire388(reg195));
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(reg174)))
        begin
          for (forvar677 = (1'h0); (forvar677 < (3'h4)); forvar677 = (forvar677 + (1'h1)))
            begin
              reg678 = (|$signed((reg190 | ((8'hb2) <<< (reg195 ?
                  wire24 : reg193)))));
              reg679 = (wire322 ?
                  ((reg199 && {reg203[(4'hb):(2'h3)], {wire169, forvar192}}) ?
                      (reg197[(5'h10):(4'hd)] ?
                          (!{wire323}) : $signed($signed(wire323))) : $signed($unsigned(wire675))) : {$unsigned(wire26)});
              reg680 <= {((!(wire323[(3'h6):(1'h1)] ?
                      (reg173 ?
                          (8'hba) : reg202) : $unsigned(forvar195))) != $signed($unsigned($unsigned(wire26))))};
              reg681 <= (~&reg177[(4'h8):(1'h1)]);
              reg682 <= (^~(^~forvar199[(2'h2):(1'h1)]));
            end
        end
      else
        begin
          for (forvar677 = (1'h0); (forvar677 < (3'h4)); forvar677 = (forvar677 + (1'h1)))
            begin
              reg678 <= $unsigned($unsigned($unsigned((reg198[(2'h2):(1'h1)] + $signed(wire324)))));
            end
          for (forvar679 = (1'h0); (forvar679 < (1'h0)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 <= ((!{forvar180, $signed($signed((8'hb2)))}) ?
                  {$unsigned($unsigned((!forvar181))),
                      $signed(($signed(reg678) ?
                          forvar181[(2'h3):(1'h0)] : (reg175 ?
                              reg202 : forvar188)))} : reg203);
              reg681 <= reg183;
            end
          reg682 <= ((reg682 | $unsigned($signed((!wire325)))) ?
              (~reg177[(5'h13):(2'h2)]) : $signed((^($unsigned((8'ha7)) != $signed(reg178)))));
        end
      reg683 <= $signed(({forvar171[(4'ha):(1'h0)]} >= ($signed((wire23 >= wire25)) ?
          (~&(~^wire675)) : (-(|wire23)))));
      for (forvar684 = (1'h0); (forvar684 < (2'h3)); forvar684 = (forvar684 + (1'h1)))
        begin
          reg685 = ($signed(reg203) ?
              (($unsigned((reg184 >= reg193)) >>> wire325) > {(8'h9f),
                  (((8'hbe) ?
                      forvar195 : reg174) - reg191)}) : (&$unsigned(($unsigned((8'ha0)) | (reg194 ?
                  wire324 : reg194)))));
          if ((~|wire325[(2'h2):(1'h1)]))
            begin
              reg686 <= (^~reg183);
              reg687 = $unsigned({(reg195[(5'h11):(5'h10)] ?
                      ("nAZdPmx4a4irKLd4Yl04" ^ reg683[(5'h12):(4'he)]) : $unsigned(reg196[(4'h8):(2'h3)]))});
            end
          else
            begin
              reg686 = ((~&(~&reg192[(2'h2):(1'h0)])) ?
                  wire325[(4'h9):(4'h9)] : $signed(wire23));
            end
          reg688 <= (reg198 ?
              wire320 : $signed($signed($unsigned((reg680 ?
                  forvar684 : (7'h40))))));
          reg689 = ($unsigned($signed({reg177, $signed((8'ha5))})) ?
              $signed({($signed(reg683) ? $unsigned(reg178) : {(8'ha4)}),
                  (^(reg184 | wire325))}) : (wire169[(4'hc):(2'h2)] && (^~$unsigned((forvar180 ?
                  forvar684 : forvar181)))));
          reg690 <= (^(!(wire24[(4'hb):(3'h4)] ^~ (&$unsigned(reg202)))));
        end
      reg691 <= (reg176[(2'h3):(1'h0)] > "41");
    end
  assign wire692 = (-reg197[(5'h11):(4'hf)]);
  always
    @(posedge clk) begin
      reg693 = $signed(reg193);
      for (forvar694 = (1'h0); (forvar694 < (2'h3)); forvar694 = (forvar694 + (1'h1)))
        begin
          reg695 = reg203;
        end
      for (forvar696 = (1'h0); (forvar696 < (1'h0)); forvar696 = (forvar696 + (1'h1)))
        begin
          reg697 = (-(((forvar180 ~^ {reg201}) ?
                  $unsigned((8'hb7)) : (~$unsigned(wire383))) ?
              wire26[(4'he):(4'he)] : (forvar187 + {(~&reg183), {reg201}})));
          for (forvar698 = (1'h0); (forvar698 < (3'h4)); forvar698 = (forvar698 + (1'h1)))
            begin
              reg699 <= (reg184 ?
                  (&reg686[(2'h3):(2'h2)]) : (reg176[(1'h1):(1'h1)] ?
                      $signed({$unsigned((8'ha2)),
                          (|reg691)}) : reg685[(1'h1):(1'h1)]));
              reg700 <= forvar195[(4'h9):(4'h8)];
              reg701 = reg192;
              reg702 <= (8'ha0);
            end
          for (forvar703 = (1'h0); (forvar703 < (2'h2)); forvar703 = (forvar703 + (1'h1)))
            begin
              reg704 <= (8'hbe);
            end
          for (forvar705 = (1'h0); (forvar705 < (1'h1)); forvar705 = (forvar705 + (1'h1)))
            begin
              reg706 = ($unsigned({(~&reg195),
                  (~|$signed(reg194))}) > $unsigned($unsigned(forvar696[(3'h7):(3'h5)])));
              reg707 = reg699[(2'h2):(1'h0)];
              reg708 = (-{(~|$signed($signed((7'h40))))});
              reg709 = (~&$unsigned({reg198,
                  (wire26[(4'hb):(2'h3)] >>> (reg182 >>> (8'hb2)))}));
              reg710 = $unsigned(((wire169 != forvar187) ^ wire320[(4'hb):(3'h6)]));
            end
        end
      if ($signed($signed(reg203[(5'h11):(2'h3)])))
        begin
          if (wire169[(3'h4):(1'h0)])
            begin
              reg711 <= (~&wire323);
            end
          else
            begin
              reg711 <= ({((reg690[(2'h3):(1'h0)] ?
                          (reg199 != wire324) : forvar199[(2'h2):(2'h2)]) ?
                      reg185 : reg178),
                  reg711} || $unsigned((~&(reg697 ^ reg690[(1'h0):(1'h0)]))));
            end
        end
      else
        begin
          for (forvar711 = (1'h0); (forvar711 < (2'h3)); forvar711 = (forvar711 + (1'h1)))
            begin
              reg712 = {reg693};
              reg713 <= (reg183[(4'h8):(3'h5)] > reg693);
              reg714 <= (reg201 | reg689[(2'h3):(1'h1)]);
              reg715 = ("PgIC4buIKFTDuJB3PwD3" ?
                  $signed((|((forvar187 ?
                      (8'h9d) : (8'h9e)) << $unsigned(wire23)))) : reg709);
              reg716 = reg195;
            end
          if (wire169)
            begin
              reg717 = $signed($signed(reg199));
              reg718 = $signed($unsigned(reg190[(4'h9):(3'h7)]));
            end
          else
            begin
              reg717 <= forvar199;
            end
          if ($signed((~|$unsigned($unsigned((~^(8'hbf)))))))
            begin
              reg719 <= (((-$signed(reg689)) ?
                      forvar188[(3'h6):(1'h0)] : (&({(8'ha0), reg709} ?
                          reg712 : {reg685}))) ?
                  $unsigned((8'ha2)) : $signed(reg711));
            end
          else
            begin
              reg719 <= forvar171;
              reg720 <= reg174[(2'h3):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar721 = (1'h0); (forvar721 < (1'h0)); forvar721 = (forvar721 + (1'h1)))
        begin
          if (reg172[(1'h1):(1'h0)])
            begin
              reg722 <= (-(+$unsigned($signed($signed(reg710)))));
            end
          else
            begin
              reg722 = $unsigned(($unsigned(((|reg176) - (!reg700))) ?
                  wire383 : reg718[(5'h14):(5'h12)]));
              reg723 <= $unsigned(((reg687 << $signed(wire324[(3'h5):(1'h0)])) ?
                  $signed(reg686[(2'h2):(1'h0)]) : wire323[(4'ha):(3'h4)]));
              reg724 <= $unsigned($signed($unsigned((&reg695))));
              reg725 = $unsigned($unsigned(((~|(reg178 & reg697)) * $unsigned(reg702[(2'h3):(2'h3)]))));
            end
          for (forvar726 = (1'h0); (forvar726 < (3'h4)); forvar726 = (forvar726 + (1'h1)))
            begin
              reg727 <= $unsigned(reg184[(1'h1):(1'h0)]);
              reg728 = reg175;
              reg729 <= ((~&$unsigned((~^$unsigned(reg681)))) ?
                  ($signed((reg679[(2'h3):(1'h1)] ?
                      {reg702,
                          reg701} : reg713[(4'h8):(4'h8)])) << $unsigned((~&$signed(reg720)))) : ($signed($unsigned((-reg711))) * reg725[(3'h6):(1'h0)]));
              reg730 = (~^(~&(~^$signed(reg687))));
              reg731 <= $signed((~&(wire323 ?
                  ((forvar180 ? forvar703 : reg715) ?
                      {reg722,
                          reg182} : reg184[(4'h9):(4'h9)]) : reg704[(1'h0):(1'h0)])));
            end
          for (forvar732 = (1'h0); (forvar732 < (2'h3)); forvar732 = (forvar732 + (1'h1)))
            begin
              reg733 = $unsigned((|reg190));
              reg734 <= ((~^$unsigned((^~(~^reg697)))) == ({(reg691 ^~ (&reg719))} ?
                  reg719 : ((^~$signed(reg711)) ?
                      $unsigned(reg707[(4'ha):(3'h5)]) : (8'hac))));
              reg735 = ({$signed(reg716)} ^~ $unsigned((("t3CiA3FU3sXqO" ?
                  $unsigned(reg175) : $signed((8'had))) > $unsigned((~&reg708)))));
              reg736 = (8'ha3);
              reg737 <= (8'ha9);
            end
          for (forvar738 = (1'h0); (forvar738 < (2'h3)); forvar738 = (forvar738 + (1'h1)))
            begin
              reg739 <= reg727[(1'h0):(1'h0)];
              reg740 <= (($unsigned($signed((reg737 ?
                  reg179 : (8'hbe)))) >> ({{reg701, forvar711},
                  $signed(reg681)} >> $signed($unsigned(reg724)))) << reg198[(3'h6):(1'h1)]);
              reg741 = (!$signed({reg723, $unsigned(reg183[(1'h1):(1'h0)])}));
              reg742 <= (^~$unsigned(forvar188));
            end
        end
      for (forvar743 = (1'h0); (forvar743 < (1'h0)); forvar743 = (forvar743 + (1'h1)))
        begin
          for (forvar744 = (1'h0); (forvar744 < (2'h3)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= $signed({(forvar199 ?
                      reg723 : $signed(reg200[(3'h7):(2'h3)]))});
            end
          reg746 <= $unsigned((reg693 + forvar732[(4'hf):(4'ha)]));
          reg747 <= $unsigned(((((8'ha6) ?
              reg725[(3'h4):(2'h2)] : (reg739 || forvar181)) >>> (~^((8'ha4) <<< reg699))) ^~ {$unsigned($signed(reg734))}));
          if (((^$signed(forvar195)) ?
              $unsigned(reg723) : $signed((!($signed((8'hba)) ?
                  forvar744 : (forvar694 ~^ (8'ha5)))))))
            begin
              reg748 <= (-$signed(($signed(reg709[(1'h1):(1'h0)]) >>> reg184)));
              reg749 = $unsigned((reg723[(4'h8):(3'h7)] | $signed(forvar192[(4'h9):(3'h6)])));
              reg750 <= ((reg725 && $unsigned((-reg198))) >= (7'h40));
            end
          else
            begin
              reg748 <= ((reg714[(2'h2):(1'h1)] ?
                      (^~(|forvar732[(1'h1):(1'h1)])) : (8'had)) ?
                  {$unsigned((+(forvar732 == reg680)))} : {(^~forvar732),
                      (&(wire692 && (reg199 ? wire675 : reg745)))});
              reg749 = reg688;
            end
          reg751 <= ((~|(reg683 ^ ("fkmkOcBNx" != ((8'hb5) != reg176)))) * wire325);
        end
    end
  assign wire752 = wire23;
  assign wire753 = "wO6IdiOrK6HZHic4C";
  assign wire754 = $signed($signed((reg191[(3'h6):(1'h0)] <= ($unsigned(reg745) ^ $unsigned(forvar721)))));
  module326 modinst756 (wire755, clk, wire675, reg178, reg749, reg714, reg734);
  assign wire757 = (7'h44);
  module385 modinst759 (.wire389(reg749), .y(wire758), .wire386(reg700), .wire390(forvar696), .wire388(wire324), .clk(clk), .wire387(reg174));
  always
    @(posedge clk) begin
      reg760 <= $signed(((-((~&forvar181) * $unsigned(reg179))) ?
          $signed({wire23[(4'h8):(3'h5)],
              "9WRknLyMJFxBS6S1"}) : (forvar696[(4'ha):(3'h5)] ?
              reg177[(4'hf):(4'hb)] : {$unsigned((8'hb8)),
                  reg192[(3'h6):(2'h2)]})));
      reg761 <= reg706;
      for (forvar762 = (1'h0); (forvar762 < (2'h2)); forvar762 = (forvar762 + (1'h1)))
        begin
          for (forvar763 = (1'h0); (forvar763 < (1'h1)); forvar763 = (forvar763 + (1'h1)))
            begin
              reg764 <= reg173;
            end
          reg765 = (8'had);
          for (forvar766 = (1'h0); (forvar766 < (2'h3)); forvar766 = (forvar766 + (1'h1)))
            begin
              reg767 <= $signed($signed($unsigned({(reg737 ? reg683 : reg731),
                  (reg693 ? reg727 : reg739)})));
              reg768 <= "u863ezskqXR2";
            end
          for (forvar769 = (1'h0); (forvar769 < (1'h1)); forvar769 = (forvar769 + (1'h1)))
            begin
              reg770 = reg724;
              reg771 <= ($signed(wire758[(4'h9):(4'h8)]) + (^$signed($signed((reg747 - wire692)))));
              reg772 <= reg722[(1'h1):(1'h0)];
            end
          reg773 <= reg729[(5'h11):(5'h10)];
        end
      reg774 = $signed(($signed((-(reg735 << reg191))) < (-(|(reg768 ?
          (8'ha8) : reg747)))));
      for (forvar775 = (1'h0); (forvar775 < (1'h1)); forvar775 = (forvar775 + (1'h1)))
        begin
          reg776 = (reg176[(3'h4):(2'h3)] ^ (reg189[(3'h5):(1'h0)] <<< ($signed({reg678}) ?
              reg701[(2'h2):(2'h2)] : (|(reg720 < reg749)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar777 = (1'h0); (forvar777 < (2'h2)); forvar777 = (forvar777 + (1'h1)))
        begin
          if ($signed(reg202))
            begin
              reg778 = $signed($unsigned($unsigned(reg178[(3'h5):(3'h5)])));
            end
          else
            begin
              reg778 <= (reg172 ?
                  {$unsigned(($signed(reg179) ?
                          $signed(reg689) : (reg681 <= (8'hb4))))} : {(&reg702)});
              reg779 = {$unsigned(reg731[(1'h0):(1'h0)])};
            end
          reg780 = reg701;
          if ((((7'h41) ?
                  ($signed($unsigned(reg771)) ?
                      $signed(reg175[(4'hb):(4'h9)]) : (^wire24)) : ($signed($unsigned((8'had))) < (7'h41))) ?
              (&$unsigned(forvar698)) : reg717))
            begin
              reg781 <= reg194[(4'h9):(3'h4)];
              reg782 <= $signed((8'ha1));
            end
          else
            begin
              reg781 <= $unsigned(reg678);
              reg782 <= ((^(((reg739 ? reg710 : wire383) ?
                  (&forvar696) : $unsigned((8'hae))) > reg723)) == $signed({reg191,
                  ("QCrie2cvthNyJdB" ? $unsigned(reg691) : $signed((8'hb8)))}));
              reg783 <= reg192[(4'hc):(1'h0)];
              reg784 = {(($unsigned($unsigned((8'hb7))) <<< $signed((~|reg202))) ?
                      wire692 : (reg680[(3'h7):(2'h3)] ~^ $unsigned(reg192)))};
              reg785 = reg740[(4'h9):(1'h1)];
            end
          for (forvar786 = (1'h0); (forvar786 < (2'h3)); forvar786 = (forvar786 + (1'h1)))
            begin
              reg787 = reg735[(3'h5):(1'h0)];
              reg788 = ((reg787 ?
                      ($unsigned((reg203 <= forvar703)) ?
                          $signed(reg747[(1'h1):(1'h0)]) : "lhqUZlR") : $unsigned(reg713[(4'h8):(2'h3)])) ?
                  ($signed((&{reg192,
                      reg686})) == reg730) : $unsigned((reg737[(1'h1):(1'h0)] ~^ ((~&reg776) ?
                      $signed(reg767) : ((8'ha3) <= reg175)))));
              reg789 = wire758;
              reg790 <= wire24;
            end
        end
      if ((8'hba))
        begin
          if (reg779)
            begin
              reg791 = ((((!reg749[(1'h0):(1'h0)]) ?
                  reg719 : {((8'ha0) ?
                          reg687 : forvar199)}) << reg779[(3'h4):(1'h0)]) != forvar777);
              reg792 <= $unsigned("rPkaPFXudww7lDGiz");
              reg793 = {(~forvar181),
                  ({(&reg776)} ?
                      $signed(($unsigned(reg737) ?
                          $signed((8'ha9)) : (forvar684 ?
                              reg689 : reg768))) : $signed(reg745[(4'hd):(4'hd)]))};
              reg794 <= (^~(~reg196[(5'h11):(3'h5)]));
            end
          else
            begin
              reg791 <= $signed(reg742[(4'h8):(3'h7)]);
              reg792 <= forvar726;
            end
          reg795 = (~&wire322);
          for (forvar796 = (1'h0); (forvar796 < (1'h1)); forvar796 = (forvar796 + (1'h1)))
            begin
              reg797 <= $unsigned("y8SchcN2SOrqqDQ");
              reg798 <= {wire383,
                  $signed(({$signed(reg687)} ?
                      $signed($unsigned(reg699)) : "h9wr2kb"))};
              reg799 <= reg794;
              reg800 <= ({$signed($signed((reg739 ? reg185 : reg789))),
                      {(8'ha8)}} ?
                  ({(^reg719[(3'h4):(2'h3)])} == (~^$unsigned(((8'ha7) ?
                      reg702 : reg190)))) : wire675);
            end
          if (($signed($unsigned($unsigned((reg706 || reg728)))) ?
              reg735 : ({$signed($signed((8'ha1))), reg183[(3'h4):(3'h4)]} ?
                  forvar766 : (8'hbc))))
            begin
              reg801 <= (reg697 ^ (reg733[(3'h5):(3'h5)] >= (8'h9c)));
              reg802 = forvar732;
            end
          else
            begin
              reg801 <= (!$signed((|$signed((&wire24)))));
              reg802 <= reg751;
              reg803 = $unsigned($unsigned((($signed((8'ha1)) ?
                  (wire753 | (8'hb2)) : reg683) ~^ $signed((reg708 & (8'h9d))))));
            end
          if ((wire324 && reg742[(3'h4):(1'h1)]))
            begin
              reg804 <= {{wire325, $signed({(reg690 ? forvar743 : reg760)})},
                  (~^reg781)};
            end
          else
            begin
              reg804 <= ($unsigned($signed((reg724 ?
                  $signed(reg715) : $signed(reg735)))) & $unsigned(({(~^reg192),
                  (forvar180 ? reg177 : (8'hac))} - reg774[(4'h9):(3'h7)])));
              reg805 <= $signed(reg782[(3'h5):(1'h0)]);
              reg806 <= (8'haf);
              reg807 <= $signed({$unsigned({reg185, forvar796}),
                  ((~^{(8'ha5)}) ^~ (~^$unsigned((8'hae))))});
              reg808 <= {reg780};
            end
        end
      else
        begin
          for (forvar791 = (1'h0); (forvar791 < (1'h0)); forvar791 = (forvar791 + (1'h1)))
            begin
              reg792 <= $unsigned((-($unsigned(((8'ha0) >> wire324)) ?
                  (~$unsigned(wire752)) : ({reg733, wire320} > ((8'hb3) ?
                      (7'h44) : reg787)))));
              reg793 = (({reg735} ^~ reg192[(4'hd):(4'h9)]) ~^ ((~^$unsigned(forvar711)) >>> {forvar762}));
              reg794 <= ($signed(((8'hbc) ?
                  reg773[(3'h7):(3'h5)] : $unsigned((wire755 < forvar786)))) == ((~|(forvar188 ?
                  $unsigned(reg781) : $unsigned(reg771))) >> (^~reg174)));
              reg795 <= reg751;
            end
        end
      if ($signed((-(+"x9EI8TEP7p0JTazy"))))
        begin
          for (forvar809 = (1'h0); (forvar809 < (2'h2)); forvar809 = (forvar809 + (1'h1)))
            begin
              reg810 <= (forvar766 < ({(~^((8'hb0) ?
                      wire692 : (8'hbc)))} >> (^~(!((8'hb0) <<< reg709)))));
              reg811 = wire169[(1'h0):(1'h0)];
            end
          for (forvar812 = (1'h0); (forvar812 < (1'h1)); forvar812 = (forvar812 + (1'h1)))
            begin
              reg813 = (reg788 ?
                  (^~"RSegO") : $signed({((~reg768) || $signed((8'hac))),
                      reg678}));
            end
          reg814 <= $unsigned((-($signed(forvar791[(5'h10):(4'h9)]) - (+$unsigned(reg749)))));
          reg815 = ($unsigned("wYdcUAnbt4wT") << $unsigned(reg176[(1'h0):(1'h0)]));
        end
      else
        begin
          for (forvar809 = (1'h0); (forvar809 < (2'h2)); forvar809 = (forvar809 + (1'h1)))
            begin
              reg810 <= ((reg751[(1'h0):(1'h0)] > wire325[(4'hb):(4'hb)]) ?
                  (((!$unsigned(forvar171)) ?
                          reg728[(2'h2):(2'h2)] : $signed({wire23})) ?
                      ($unsigned((reg781 ?
                          wire26 : reg701)) >> (+reg173)) : ($unsigned("G6BvONLmoRe4dwPbA") & $unsigned((|reg185)))) : (~&(+$unsigned($unsigned(reg790)))));
              reg811 <= $unsigned("Qd");
              reg812 = (&$unsigned($unsigned($unsigned((~|reg761)))));
            end
          reg813 <= $signed($signed({reg193}));
          reg814 <= (~^{({reg706[(1'h0):(1'h0)]} << $unsigned(reg733))});
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module385
#( parameter param673 = (((((~&(8'h9c)) <<< ((8'hba) * (8'ha2))) ? (((8'hb0) * (8'hb7)) <<< ((8'ha1) ? (7'h42) : (7'h43))) : (~|((8'hac) ? (8'hb6) : (8'hb6)))) > ((((8'hb4) ? (8'hb7) : (7'h40)) ? ((7'h40) != (7'h41)) : (8'hb9)) & (~((8'hbd) ? (8'ha6) : (8'hac))))) ? (^~((((8'hac) ? (8'ha3) : (8'hb6)) && ((7'h40) <<< (8'hbd))) ? (((8'hb7) >= (8'hbe)) ^ ((8'ha0) > (8'ha6))) : (^(^~(8'ha5))))) : ({(+(^~(8'ha8)))} > {((~(8'ha7)) ? ((8'hb5) > (8'ha5)) : (^(8'hb6)))}))
, parameter param674 = (((8'hb5) <= {(^~(param673 <= param673)), (^~(8'ha4))}) <<< (({(param673 ? (8'h9c) : (8'hb9))} ? ((8'hbf) < param673) : ((~^param673) ? (^~param673) : (~&(8'haa)))) ? {{param673, (param673 ? param673 : param673)}} : (~(^(!param673))))) )
(y, clk, wire390, wire389, wire388, wire387, wire386);
  output wire [(32'hd40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire390;
  input wire [(5'h14):(1'h0)] wire389;
  input wire signed [(5'h15):(1'h0)] wire388;
  input wire signed [(4'he):(1'h0)] wire387;
  input wire signed [(4'hb):(1'h0)] wire386;
  reg signed [(2'h3):(1'h0)] reg672 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg671 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg669 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg667 = (1'h0);
  reg [(4'hc):(1'h0)] forvar666 = (1'h0);
  reg [(5'h15):(1'h0)] reg665 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg664 = (1'h0);
  reg [(5'h12):(1'h0)] reg663 = (1'h0);
  reg [(3'h6):(1'h0)] reg662 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg661 = (1'h0);
  reg [(4'h8):(1'h0)] reg660 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg659 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar658 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg657 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg656 = (1'h0);
  reg [(4'hc):(1'h0)] reg655 = (1'h0);
  reg [(4'hc):(1'h0)] reg654 = (1'h0);
  reg [(4'hb):(1'h0)] forvar653 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar652 = (1'h0);
  reg [(5'h11):(1'h0)] reg651 = (1'h0);
  reg [(2'h2):(1'h0)] reg650 = (1'h0);
  reg [(4'ha):(1'h0)] reg649 = (1'h0);
  reg [(3'h5):(1'h0)] reg648 = (1'h0);
  reg [(4'he):(1'h0)] reg647 = (1'h0);
  reg [(5'h11):(1'h0)] reg646 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg645 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg644 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg643 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg642 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar641 = (1'h0);
  reg [(4'h9):(1'h0)] reg640 = (1'h0);
  reg [(4'hf):(1'h0)] reg639 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg638 = (1'h0);
  reg [(4'hf):(1'h0)] reg637 = (1'h0);
  reg [(5'h11):(1'h0)] reg636 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar634 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg632 = (1'h0);
  reg [(4'he):(1'h0)] reg631 = (1'h0);
  reg [(3'h4):(1'h0)] forvar630 = (1'h0);
  reg signed [(4'he):(1'h0)] reg629 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar628 = (1'h0);
  reg [(2'h3):(1'h0)] reg627 = (1'h0);
  reg [(5'h14):(1'h0)] reg626 = (1'h0);
  reg signed [(4'he):(1'h0)] reg625 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg624 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg623 = (1'h0);
  reg [(3'h5):(1'h0)] forvar622 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire621;
  reg signed [(4'hb):(1'h0)] reg620 = (1'h0);
  reg [(3'h5):(1'h0)] reg619 = (1'h0);
  reg [(4'he):(1'h0)] reg618 = (1'h0);
  reg [(5'h12):(1'h0)] reg617 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg616 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg615 = (1'h0);
  reg [(4'he):(1'h0)] forvar614 = (1'h0);
  reg [(4'ha):(1'h0)] forvar613 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg612 = (1'h0);
  reg [(4'h8):(1'h0)] reg611 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar609 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg608 = (1'h0);
  reg [(4'h8):(1'h0)] reg607 = (1'h0);
  reg signed [(4'he):(1'h0)] reg606 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg605 = (1'h0);
  reg [(5'h13):(1'h0)] forvar604 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg603 = (1'h0);
  reg [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(3'h6):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar600 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg599 = (1'h0);
  reg [(5'h11):(1'h0)] reg598 = (1'h0);
  reg [(3'h7):(1'h0)] reg597 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg595 = (1'h0);
  reg [(4'he):(1'h0)] reg594 = (1'h0);
  reg [(5'h15):(1'h0)] forvar593 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg592 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg591 = (1'h0);
  reg [(4'ha):(1'h0)] reg590 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg588 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar587 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg586 = (1'h0);
  reg [(3'h7):(1'h0)] reg585 = (1'h0);
  reg [(3'h7):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg583 = (1'h0);
  reg [(4'he):(1'h0)] reg582 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg581 = (1'h0);
  reg [(5'h14):(1'h0)] reg580 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar579 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire578;
  wire signed [(4'h9):(1'h0)] wire577;
  reg signed [(4'he):(1'h0)] reg576 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg573 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar572 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg571 = (1'h0);
  reg [(5'h13):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg569 = (1'h0);
  reg [(4'h8):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar567 = (1'h0);
  reg [(4'hf):(1'h0)] forvar566 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar560 = (1'h0);
  reg [(5'h15):(1'h0)] reg565 = (1'h0);
  reg [(5'h11):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg563 = (1'h0);
  reg [(4'hd):(1'h0)] reg562 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg561 = (1'h0);
  reg [(5'h13):(1'h0)] reg560 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg559 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar558 = (1'h0);
  reg [(2'h3):(1'h0)] reg557 = (1'h0);
  reg [(4'hc):(1'h0)] reg556 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg555 = (1'h0);
  reg [(5'h14):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg552 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg550 = (1'h0);
  reg [(5'h11):(1'h0)] forvar549 = (1'h0);
  reg [(3'h6):(1'h0)] reg548 = (1'h0);
  reg [(5'h13):(1'h0)] reg547 = (1'h0);
  reg [(5'h12):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg543 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar542 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg541 = (1'h0);
  reg [(5'h13):(1'h0)] reg540 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg539 = (1'h0);
  reg [(3'h6):(1'h0)] reg538 = (1'h0);
  reg [(5'h11):(1'h0)] forvar537 = (1'h0);
  reg [(3'h7):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar533 = (1'h0);
  reg [(2'h2):(1'h0)] forvar529 = (1'h0);
  reg [(5'h13):(1'h0)] reg524 = (1'h0);
  reg [(4'he):(1'h0)] reg535 = (1'h0);
  reg [(3'h5):(1'h0)] reg534 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg533 = (1'h0);
  reg [(5'h12):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg530 = (1'h0);
  reg [(3'h5):(1'h0)] reg529 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg528 = (1'h0);
  reg [(5'h13):(1'h0)] reg527 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg526 = (1'h0);
  reg [(4'he):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar524 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg523 = (1'h0);
  reg [(2'h3):(1'h0)] reg522 = (1'h0);
  reg [(4'hc):(1'h0)] reg521 = (1'h0);
  reg signed [(4'he):(1'h0)] reg520 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg519 = (1'h0);
  reg [(3'h7):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg517 = (1'h0);
  reg signed [(4'he):(1'h0)] reg516 = (1'h0);
  reg [(2'h2):(1'h0)] reg515 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar514 = (1'h0);
  reg signed [(4'he):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar512 = (1'h0);
  reg [(4'hb):(1'h0)] forvar511 = (1'h0);
  reg [(3'h5):(1'h0)] reg510 = (1'h0);
  reg [(5'h12):(1'h0)] reg509 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar507 = (1'h0);
  reg [(5'h12):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar503 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar502 = (1'h0);
  wire signed [(4'he):(1'h0)] wire501;
  wire signed [(5'h14):(1'h0)] wire500;
  wire [(5'h13):(1'h0)] wire499;
  reg signed [(4'h9):(1'h0)] reg498 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg497 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg496 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar495 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg494 = (1'h0);
  reg [(5'h13):(1'h0)] forvar493 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg491 = (1'h0);
  reg [(5'h10):(1'h0)] reg490 = (1'h0);
  reg [(5'h15):(1'h0)] reg489 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar488 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg486 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg485 = (1'h0);
  reg [(3'h6):(1'h0)] reg484 = (1'h0);
  reg [(4'hb):(1'h0)] reg483 = (1'h0);
  reg [(4'hd):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg480 = (1'h0);
  reg [(5'h11):(1'h0)] reg479 = (1'h0);
  reg [(4'h8):(1'h0)] forvar478 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar477 = (1'h0);
  reg [(5'h11):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg [(4'hd):(1'h0)] reg474 = (1'h0);
  reg [(3'h5):(1'h0)] reg473 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg472 = (1'h0);
  reg [(4'hd):(1'h0)] forvar471 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg470 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg469 = (1'h0);
  reg [(4'h9):(1'h0)] reg468 = (1'h0);
  reg [(5'h11):(1'h0)] reg467 = (1'h0);
  reg [(3'h5):(1'h0)] forvar466 = (1'h0);
  reg [(3'h7):(1'h0)] reg465 = (1'h0);
  reg [(5'h11):(1'h0)] reg464 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg463 = (1'h0);
  reg [(5'h12):(1'h0)] reg462 = (1'h0);
  reg [(4'hb):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar460 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg459 = (1'h0);
  reg [(4'ha):(1'h0)] reg458 = (1'h0);
  reg [(5'h12):(1'h0)] forvar457 = (1'h0);
  reg [(4'he):(1'h0)] reg456 = (1'h0);
  reg [(3'h5):(1'h0)] reg455 = (1'h0);
  reg [(4'hd):(1'h0)] reg454 = (1'h0);
  reg [(5'h10):(1'h0)] reg453 = (1'h0);
  reg [(5'h12):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar451 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg450 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar449 = (1'h0);
  reg [(4'h8):(1'h0)] reg448 = (1'h0);
  reg [(3'h7):(1'h0)] forvar447 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar446 = (1'h0);
  reg [(4'hc):(1'h0)] reg441 = (1'h0);
  reg [(4'h8):(1'h0)] forvar438 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg437 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg433 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar432 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar429 = (1'h0);
  reg [(4'hf):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg445 = (1'h0);
  reg [(5'h15):(1'h0)] reg444 = (1'h0);
  reg [(4'h9):(1'h0)] reg443 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg442 = (1'h0);
  reg [(5'h15):(1'h0)] forvar441 = (1'h0);
  reg [(4'ha):(1'h0)] reg440 = (1'h0);
  reg [(2'h3):(1'h0)] reg439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg438 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar437 = (1'h0);
  reg [(4'he):(1'h0)] reg436 = (1'h0);
  reg [(4'hc):(1'h0)] reg435 = (1'h0);
  reg [(4'hf):(1'h0)] reg434 = (1'h0);
  reg [(4'hc):(1'h0)] forvar433 = (1'h0);
  reg [(2'h3):(1'h0)] reg432 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg430 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg429 = (1'h0);
  reg [(2'h2):(1'h0)] forvar428 = (1'h0);
  reg [(4'hc):(1'h0)] reg427 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg426 = (1'h0);
  reg [(5'h15):(1'h0)] reg425 = (1'h0);
  reg [(5'h14):(1'h0)] reg424 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg423 = (1'h0);
  reg signed [(4'he):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg419 = (1'h0);
  reg [(5'h12):(1'h0)] forvar418 = (1'h0);
  reg [(4'hb):(1'h0)] reg417 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg416 = (1'h0);
  reg [(5'h10):(1'h0)] reg415 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar412 = (1'h0);
  reg [(5'h13):(1'h0)] reg411 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg410 = (1'h0);
  reg signed [(4'he):(1'h0)] reg409 = (1'h0);
  reg [(5'h13):(1'h0)] reg408 = (1'h0);
  reg [(4'h8):(1'h0)] forvar407 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar406 = (1'h0);
  reg [(4'h8):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg404 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire403;
  reg [(4'h8):(1'h0)] reg402 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg393 = (1'h0);
  reg signed [(4'he):(1'h0)] reg401 = (1'h0);
  reg [(5'h15):(1'h0)] reg400 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg399 = (1'h0);
  reg [(4'hb):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg397 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg395 = (1'h0);
  reg [(4'hc):(1'h0)] reg394 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar393 = (1'h0);
  reg [(3'h7):(1'h0)] reg392 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire391;
  assign y = {reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 forvar666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 forvar658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 forvar653,
                 forvar652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 forvar641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 forvar634,
                 reg633,
                 reg632,
                 reg631,
                 forvar630,
                 reg629,
                 forvar628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 forvar622,
                 wire621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 forvar614,
                 forvar613,
                 reg612,
                 reg611,
                 reg610,
                 forvar609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 forvar604,
                 reg603,
                 reg602,
                 reg601,
                 forvar600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 forvar593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 forvar587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 wire578,
                 wire577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 forvar572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 forvar567,
                 forvar566,
                 forvar560,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 forvar558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 forvar549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 forvar542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 forvar537,
                 reg536,
                 forvar533,
                 forvar529,
                 reg524,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 forvar524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 forvar512,
                 forvar511,
                 reg510,
                 reg509,
                 reg508,
                 forvar507,
                 reg506,
                 reg505,
                 reg504,
                 forvar503,
                 forvar502,
                 wire501,
                 wire500,
                 wire499,
                 reg498,
                 reg497,
                 reg496,
                 forvar495,
                 reg494,
                 forvar493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 forvar488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 forvar478,
                 forvar477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 forvar471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 forvar466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 forvar460,
                 reg459,
                 reg458,
                 forvar457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 forvar451,
                 reg450,
                 forvar449,
                 reg448,
                 forvar447,
                 forvar446,
                 reg441,
                 forvar438,
                 reg437,
                 reg433,
                 forvar432,
                 forvar429,
                 reg428,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 forvar441,
                 reg440,
                 reg439,
                 reg438,
                 forvar437,
                 reg436,
                 reg435,
                 reg434,
                 forvar433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 forvar428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 forvar418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 forvar412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 forvar406,
                 reg405,
                 reg404,
                 wire403,
                 reg402,
                 reg393,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 reg392,
                 wire391,
                 (1'h0)};
  assign wire391 = {wire388[(5'h14):(5'h10)]};
  always
    @(posedge clk) begin
      reg392 = wire387[(4'hc):(4'ha)];
      if (((&(reg392[(3'h7):(3'h7)] ?
              ({wire390} ?
                  (wire391 >= wire388) : (wire388 == (8'ha5))) : $unsigned(wire386))) ?
          $signed((~&((!wire386) != wire386))) : $signed($signed($unsigned((wire387 ?
              reg392 : (8'hb0)))))))
        begin
          for (forvar393 = (1'h0); (forvar393 < (2'h3)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= $signed(wire390);
              reg395 = reg394[(2'h3):(1'h0)];
              reg396 <= wire390[(3'h7):(3'h4)];
            end
          if ($signed($signed(wire391)))
            begin
              reg397 <= forvar393[(1'h0):(1'h0)];
              reg398 <= wire389;
              reg399 = $unsigned((~($signed((reg394 ? wire390 : reg397)) ?
                  (|$unsigned(reg395)) : (wire388 ?
                      ((8'ha4) <<< wire389) : (+wire391)))));
              reg400 = (+wire389[(4'hf):(2'h3)]);
              reg401 <= reg392[(3'h4):(2'h3)];
            end
          else
            begin
              reg397 = (~^(8'hb2));
              reg398 <= $unsigned(reg392);
              reg399 = (~^wire387);
              reg400 <= $signed(wire388);
            end
        end
      else
        begin
          if (wire390[(3'h7):(2'h3)])
            begin
              reg393 <= $signed(($unsigned($unsigned({reg395,
                  wire389})) >> reg397[(2'h2):(1'h1)]));
              reg394 = (((^$unsigned($unsigned(wire386))) ?
                      ($unsigned((+forvar393)) ?
                          $signed({wire386}) : {(reg399 ?
                                  (8'h9f) : (8'hae))}) : ((+$signed(reg398)) ^~ ((8'h9f) >> (reg394 ?
                          wire386 : reg395)))) ?
                  $unsigned($unsigned((8'h9c))) : reg394);
              reg395 <= (~(&$signed(((-reg392) << $unsigned(reg397)))));
              reg396 = $signed($signed((({(8'hb4)} <= $signed(wire386)) ?
                  reg393[(3'h5):(1'h0)] : "D")));
              reg397 = reg398;
            end
          else
            begin
              reg393 <= (($unsigned(wire389) ?
                      (reg394[(4'hb):(2'h3)] | $unsigned((~reg398))) : (!($signed(reg398) ?
                          (wire386 > reg397) : $unsigned(reg393)))) ?
                  ({wire386[(4'h8):(3'h7)],
                          {$unsigned(reg399), (wire386 + wire386)}} ?
                      $signed($unsigned((reg395 ?
                          reg393 : (8'ha9)))) : (((reg392 ?
                              wire390 : reg393) || (8'ha0)) ?
                          $unsigned((wire389 ? wire389 : (8'hbb))) : ((wire387 ?
                              wire388 : reg401) >>> $signed(reg395)))) : $unsigned((&(-reg394[(4'hb):(3'h6)]))));
            end
          reg398 = $signed($unsigned(wire387[(2'h3):(1'h1)]));
          reg399 <= ((8'hbe) != (reg396 ?
              ($unsigned(reg393[(1'h0):(1'h0)]) < ($unsigned((7'h43)) ^~ (!wire386))) : (((wire387 == (8'h9f)) ?
                      (&(8'ha6)) : wire390) ?
                  {forvar393[(4'h9):(3'h7)],
                      $signed(reg399)} : reg396[(2'h2):(1'h1)])));
        end
      reg402 = reg395;
    end
  assign wire403 = ($unsigned((reg400 >= reg393[(3'h4):(1'h0)])) + {{{$unsigned(wire389),
                               (-wire390)}}});
  always
    @(posedge clk) begin
      reg404 = wire388[(1'h1):(1'h0)];
      reg405 = ((^(wire386 ?
          ((wire389 ?
              wire390 : wire390) < $unsigned(reg402)) : $signed((reg393 == reg396)))) >>> (~($unsigned((reg398 + wire403)) ?
          reg398[(4'h9):(4'h9)] : ($unsigned((8'ha7)) ?
              (reg402 ? (8'ha6) : (8'had)) : (reg400 ^~ reg396)))));
      for (forvar406 = (1'h0); (forvar406 < (3'h4)); forvar406 = (forvar406 + (1'h1)))
        begin
          for (forvar407 = (1'h0); (forvar407 < (1'h1)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 = (~^$signed($signed(((^~forvar406) + (|wire386)))));
              reg409 <= (^~{({(reg399 > reg408)} ?
                      $unsigned((reg396 ? reg405 : wire388)) : (|(+(7'h42))))});
              reg410 = $signed(($unsigned((forvar406[(2'h3):(1'h0)] >> $signed(reg409))) || (~&$signed(reg396[(4'h9):(3'h4)]))));
              reg411 <= forvar407[(1'h0):(1'h0)];
            end
          for (forvar412 = (1'h0); (forvar412 < (1'h1)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 = $signed($unsigned(wire389[(1'h0):(1'h0)]));
              reg414 = $unsigned(wire403);
              reg415 <= ((~$signed(({reg393, wire391} ?
                  ((8'had) ? (8'hb3) : wire389) : {reg399}))) ^~ (reg402 ?
                  $signed(reg394[(1'h0):(1'h0)]) : ($unsigned((reg414 ?
                      reg398 : reg414)) & (forvar393 <<< $signed(reg394)))));
              reg416 <= $signed($signed($unsigned(reg399[(3'h7):(1'h1)])));
              reg417 <= (&(reg410[(2'h2):(2'h2)] && $signed(reg416)));
            end
          for (forvar418 = (1'h0); (forvar418 < (2'h3)); forvar418 = (forvar418 + (1'h1)))
            begin
              reg419 <= {((reg400[(5'h14):(2'h3)] ?
                      "t6JArV" : ((~&forvar406) + {reg404,
                          forvar406})) || (reg397[(2'h2):(1'h0)] <<< ($signed(reg415) ?
                      wire389 : reg395[(2'h2):(1'h1)])))};
              reg420 = {$signed($signed((reg401 + forvar418[(1'h1):(1'h1)]))),
                  reg402[(2'h3):(1'h1)]};
              reg421 <= $unsigned(wire403[(4'hb):(3'h6)]);
              reg422 = $signed(reg411[(4'hc):(3'h7)]);
              reg423 = "";
            end
          reg424 = reg422;
          if ((reg394[(4'h9):(2'h2)] ?
              {$unsigned((reg393[(3'h5):(3'h4)] ?
                      ((8'ha7) == wire389) : (~&reg399))),
                  {""}} : (reg414[(2'h2):(1'h0)] - (wire403[(3'h4):(2'h2)] ?
                  $signed((reg395 ? reg415 : (8'ha1))) : ((forvar412 ?
                          reg423 : reg416) ?
                      $signed(reg402) : (reg416 ~^ reg398))))))
            begin
              reg425 = reg392;
              reg426 = ($unsigned($unsigned((!(reg398 ^~ wire389)))) ?
                  (^(((reg411 <<< reg417) ~^ (!reg414)) ?
                      ((+forvar412) ?
                          reg421 : wire389[(3'h7):(2'h2)]) : (~&(reg416 == reg411)))) : $unsigned((7'h41)));
            end
          else
            begin
              reg425 = $unsigned(((~{{wire390,
                      reg416}}) - ("Dtp" != $signed((|reg417)))));
              reg426 = (~&(+(forvar418 ?
                  $signed(reg394[(3'h5):(1'h1)]) : $unsigned((~&forvar412)))));
              reg427 <= (wire386 ?
                  (~&((!{forvar407,
                      reg392}) && $signed(reg419[(4'ha):(3'h4)]))) : $unsigned(reg393[(3'h5):(1'h1)]));
            end
        end
      if (wire391[(3'h4):(3'h4)])
        begin
          for (forvar428 = (1'h0); (forvar428 < (2'h3)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 <= "GEqLvrvcTGbXu5h7y0oa";
              reg430 <= reg414;
              reg431 <= (wire388 < $unsigned($unsigned(reg399[(2'h2):(1'h1)])));
              reg432 = ($signed(reg420) ?
                  $signed(((&(reg400 & reg411)) | (+(reg425 || wire389)))) : ({(reg427[(4'h9):(1'h0)] != (~^reg417)),
                      wire387[(4'h9):(3'h4)]} >= reg392[(1'h1):(1'h0)]));
            end
          for (forvar433 = (1'h0); (forvar433 < (1'h0)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= (^(~reg421[(1'h0):(1'h0)]));
              reg435 = reg434[(4'h9):(3'h6)];
              reg436 <= $unsigned({$unsigned($signed((reg430 ?
                      reg417 : reg421)))});
            end
          for (forvar437 = (1'h0); (forvar437 < (1'h1)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= $signed((($signed(reg436) ?
                  ((-reg436) == $signed((8'had))) : forvar418) - $unsigned(wire403[(3'h4):(1'h1)])));
              reg439 = $unsigned((forvar406[(4'h8):(3'h6)] || (wire388[(4'hc):(1'h1)] ?
                  (&reg414) : (~^(reg420 ? reg429 : reg426)))));
              reg440 <= ((^(^~{$unsigned(wire391),
                  (-reg410)})) << $unsigned(("O02hqzmZQGcbMt3t" ^ (reg415 - reg416))));
            end
          for (forvar441 = (1'h0); (forvar441 < (3'h4)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 = {$unsigned((!((forvar393 << wire389) ?
                      (-reg417) : reg430)))};
              reg443 = {(forvar428 | $signed(((|(8'hb0)) - forvar412))),
                  (~&(reg430 != reg422[(4'ha):(4'h9)]))};
              reg444 = (({$signed((^forvar418))} << (+$signed((8'h9c)))) ?
                  forvar407 : reg401[(3'h4):(2'h3)]);
            end
          reg445 <= (reg408[(3'h5):(2'h2)] ?
              forvar441 : $signed("3LMXIbMpVxIW"));
        end
      else
        begin
          reg428 <= ($unsigned(reg438) << $signed(reg436));
          for (forvar429 = (1'h0); (forvar429 < (1'h1)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 = reg392;
              reg431 <= $unsigned($unsigned($unsigned(reg428[(2'h2):(2'h2)])));
            end
          for (forvar432 = (1'h0); (forvar432 < (2'h2)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= (|({{$unsigned(reg420),
                      $unsigned(reg429)}} <= (reg422 <<< $unsigned({wire390,
                  reg399}))));
              reg434 <= reg413;
              reg435 <= "lfye5D";
              reg436 = {reg410[(2'h3):(1'h1)], (|reg416)};
              reg437 <= ({(((reg410 ? wire391 : reg440) >>> $signed(reg427)) ?
                      {$signed(wire386),
                          {forvar428, reg402}} : ($unsigned(reg431) ?
                          (reg433 != reg421) : $signed(forvar433))),
                  ((&{reg405}) | forvar437[(1'h0):(1'h0)])} || $signed($unsigned(forvar441)));
            end
          for (forvar438 = (1'h0); (forvar438 < (3'h4)); forvar438 = (forvar438 + (1'h1)))
            begin
              reg439 = $signed((~^($signed(reg445[(4'hc):(4'ha)]) ?
                  $unsigned($unsigned(reg424)) : reg400)));
              reg440 <= reg433[(1'h1):(1'h0)];
            end
          reg441 <= {reg416[(3'h4):(1'h1)]};
        end
    end
  always
    @(posedge clk) begin
      for (forvar446 = (1'h0); (forvar446 < (2'h2)); forvar446 = (forvar446 + (1'h1)))
        begin
          for (forvar447 = (1'h0); (forvar447 < (1'h1)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 <= wire388[(1'h1):(1'h0)];
            end
          for (forvar449 = (1'h0); (forvar449 < (3'h4)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 <= forvar428;
            end
          for (forvar451 = (1'h0); (forvar451 < (1'h1)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 <= ({(!(+(|forvar438)))} * $signed("gErq"));
              reg453 = ((reg424 & {((~|reg444) ?
                          (+reg392) : (wire389 >>> (8'hbe))),
                      (reg424[(4'hd):(4'hd)] ?
                          $signed(wire390) : (reg450 ? (8'ha0) : reg429))}) ?
                  ($unsigned($unsigned((wire389 - reg405))) <<< (($signed(reg452) ^ (~|reg450)) < $unsigned((^~reg415)))) : reg438);
              reg454 <= reg410[(1'h0):(1'h0)];
              reg455 <= $signed(reg413);
              reg456 <= reg395[(3'h5):(1'h0)];
            end
        end
      for (forvar457 = (1'h0); (forvar457 < (1'h0)); forvar457 = (forvar457 + (1'h1)))
        begin
          reg458 <= ($signed($unsigned(reg398[(3'h6):(3'h4)])) ?
              reg435[(4'h9):(1'h0)] : {(-reg395[(3'h4):(2'h2)]),
                  $signed((8'h9f))});
          reg459 <= (&(reg427[(3'h7):(1'h1)] ?
              $signed($unsigned(reg404[(3'h5):(3'h4)])) : $unsigned(($signed(reg414) < $signed(reg435)))));
          for (forvar460 = (1'h0); (forvar460 < (2'h3)); forvar460 = (forvar460 + (1'h1)))
            begin
              reg461 = (reg417[(1'h1):(1'h0)] ^ (^($signed(reg448[(2'h2):(2'h2)]) ?
                  $signed({reg410}) : (wire391[(2'h2):(2'h2)] >= reg443))));
              reg462 <= ({reg438[(2'h2):(1'h1)]} ? reg424 : (&wire391));
              reg463 <= forvar433[(4'h8):(4'h8)];
              reg464 <= ($signed((^~$unsigned($signed(reg409)))) ?
                  (-(8'hb3)) : forvar460);
              reg465 <= (reg421 >> $unsigned((~((forvar446 ?
                      forvar457 : forvar429) ?
                  reg435 : (+forvar393)))));
            end
        end
      for (forvar466 = (1'h0); (forvar466 < (2'h3)); forvar466 = (forvar466 + (1'h1)))
        begin
          if ((~^($unsigned(((reg453 >= reg399) ?
              $unsigned(reg397) : {reg420, reg444})) <= reg459[(1'h1):(1'h1)])))
            begin
              reg467 = $signed($unsigned($unsigned(reg458)));
              reg468 = ($unsigned($signed((reg435 ^ $unsigned((8'haf))))) + ((-forvar407) <= forvar437));
              reg469 <= (8'ha1);
              reg470 = (~&forvar451);
            end
          else
            begin
              reg467 <= ((!($signed(((8'hbc) ? reg459 : forvar449)) ?
                      reg439[(2'h3):(1'h1)] : $unsigned((^~reg394)))) ?
                  "t" : $unsigned((("wXwunocc" >> {reg431}) != (reg420[(3'h7):(1'h0)] ?
                      $signed(wire390) : $unsigned(reg435)))));
              reg468 <= ((($signed(reg393) ?
                  reg440[(4'ha):(3'h4)] : {reg402}) <<< $signed($signed("7"))) <= forvar432[(1'h0):(1'h0)]);
              reg469 = (8'ha1);
              reg470 <= $signed($unsigned({reg465}));
            end
          for (forvar471 = (1'h0); (forvar471 < (3'h4)); forvar471 = (forvar471 + (1'h1)))
            begin
              reg472 <= (-(~|(~&$signed($unsigned(reg404)))));
              reg473 = reg445[(5'h13):(3'h6)];
              reg474 <= (reg396 ^~ $unsigned({$unsigned("XPVNRB"),
                  reg411[(1'h1):(1'h1)]}));
              reg475 <= $unsigned(forvar432[(3'h5):(2'h3)]);
              reg476 <= $unsigned({wire390});
            end
        end
      for (forvar477 = (1'h0); (forvar477 < (2'h3)); forvar477 = (forvar477 + (1'h1)))
        begin
          for (forvar478 = (1'h0); (forvar478 < (1'h0)); forvar478 = (forvar478 + (1'h1)))
            begin
              reg479 = (($unsigned(forvar451[(1'h1):(1'h1)]) < ($unsigned(reg422[(3'h6):(2'h3)]) >> forvar457)) >> $unsigned(wire390));
              reg480 <= reg424;
              reg481 = (reg444 >= (7'h40));
              reg482 = reg463[(4'h8):(2'h3)];
              reg483 = (+((~^((-reg431) ?
                      reg440[(4'h8):(3'h5)] : $signed((8'hb7)))) ?
                  (~(^~reg429[(1'h1):(1'h0)])) : (~|((forvar393 < forvar418) ?
                      (wire390 > reg458) : {forvar447}))));
            end
        end
      if ({(~forvar393[(3'h6):(3'h5)]), wire389})
        begin
          if ($unsigned("i1hnmOKkcgYYG"))
            begin
              reg484 <= reg392;
              reg485 = ({$signed(reg474)} ?
                  (reg427[(3'h7):(2'h2)] ?
                      reg397[(3'h4):(2'h2)] : (((forvar471 | wire390) ?
                              $unsigned(reg396) : $unsigned(forvar429)) ?
                          reg404 : (reg484[(3'h5):(3'h4)] ^~ reg437))) : forvar451);
            end
          else
            begin
              reg484 <= (~|(8'h9c));
              reg485 = reg399[(4'h8):(3'h6)];
              reg486 <= ({(reg408 ?
                      (reg401 << reg443[(1'h1):(1'h1)]) : (8'ha2))} * (+$unsigned((~$unsigned(forvar428)))));
            end
        end
      else
        begin
          if ($signed((-reg482)))
            begin
              reg484 = (reg422 ? reg455 : reg483);
              reg485 = (((!(&reg436)) ?
                  (reg469 ?
                      ($signed(forvar457) ?
                          (^~reg432) : $unsigned(wire403)) : reg428) : $signed(((~reg484) ?
                      (^(8'hb6)) : (wire390 >= (8'hac))))) && reg436);
            end
          else
            begin
              reg484 <= $unsigned(reg474);
              reg485 <= $signed(reg405[(4'h8):(1'h0)]);
              reg486 <= $signed((reg414 ?
                  $unsigned(((-reg411) ?
                      $unsigned((8'hb7)) : (forvar429 | forvar432))) : (((reg464 ?
                      reg442 : reg463) - (forvar429 ^~ (8'ha5))) <= (reg444 <= (reg437 >= reg441)))));
              reg487 <= ($signed(reg419) <<< forvar407[(3'h7):(3'h4)]);
            end
          for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
            begin
              reg489 = forvar407;
              reg490 = $signed(((reg448[(1'h0):(1'h0)] ?
                  reg437[(5'h12):(3'h4)] : reg486) >= wire390[(3'h4):(2'h2)]));
              reg491 = reg490[(4'ha):(4'h9)];
            end
          reg492 = {($signed(reg432) ?
                  {reg405[(3'h6):(2'h3)]} : (^~{"KoDXtead8OnXrmUAaVXD",
                      (reg413 ? reg464 : (8'h9e))})),
              reg489};
          for (forvar493 = (1'h0); (forvar493 < (2'h3)); forvar493 = (forvar493 + (1'h1)))
            begin
              reg494 <= "A55C0S";
            end
          for (forvar495 = (1'h0); (forvar495 < (2'h3)); forvar495 = (forvar495 + (1'h1)))
            begin
              reg496 = $unsigned(((((reg442 >= forvar471) >= (^(8'hb4))) ?
                      (+$unsigned(reg400)) : (+reg435)) ?
                  (forvar441 ?
                      (|$signed(reg420)) : $unsigned(reg415)) : reg395[(3'h5):(3'h4)]));
              reg497 <= reg395[(4'hd):(2'h2)];
              reg498 <= wire386[(1'h1):(1'h0)];
            end
        end
    end
  assign wire499 = {((($unsigned(reg422) != reg404) ?
                           ($unsigned(reg448) ?
                               forvar438[(4'h8):(4'h8)] : reg486[(4'h9):(1'h1)]) : $signed($signed(reg419))) <= $signed($signed($unsigned(reg464)))),
                       ((8'h9c) ?
                           (^$signed((-forvar446))) : reg408[(1'h0):(1'h0)])};
  assign wire500 = (({reg484} || $unsigned($unsigned($signed((7'h40))))) + forvar437);
  assign wire501 = (reg409 < forvar447[(3'h5):(2'h3)]);
  always
    @(posedge clk) begin
      for (forvar502 = (1'h0); (forvar502 < (1'h1)); forvar502 = (forvar502 + (1'h1)))
        begin
          for (forvar503 = (1'h0); (forvar503 < (1'h0)); forvar503 = (forvar503 + (1'h1)))
            begin
              reg504 = (|$unsigned((|$signed($signed((8'ha9))))));
              reg505 <= $unsigned(reg459[(2'h2):(1'h1)]);
            end
          reg506 <= (($unsigned({reg423[(2'h2):(2'h2)],
                  ((8'hbb) ? reg427 : (7'h41))}) ?
              (reg445[(4'ha):(3'h4)] || $signed($unsigned((8'h9f)))) : reg399[(4'h8):(1'h1)]) + reg486);
          for (forvar507 = (1'h0); (forvar507 < (1'h1)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 <= "ItmfiK";
            end
          reg509 = reg425[(3'h4):(2'h3)];
        end
      reg510 <= ((~^(+forvar451)) >>> $signed({reg455[(2'h2):(1'h0)],
          ((reg509 ? reg455 : reg467) ? (^reg448) : forvar471)}));
      for (forvar511 = (1'h0); (forvar511 < (3'h4)); forvar511 = (forvar511 + (1'h1)))
        begin
          for (forvar512 = (1'h0); (forvar512 < (2'h3)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 <= reg435[(4'h8):(1'h1)];
            end
          for (forvar514 = (1'h0); (forvar514 < (3'h4)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 <= "xVgvDSauC8fE6YBzh";
              reg516 <= $unsigned((reg422 <= {(~&reg422),
                  ({(8'hbd), reg504} ?
                      {reg443, wire390} : forvar432[(3'h4):(2'h3)])}));
              reg517 <= $signed((reg491 ?
                  reg416[(1'h0):(1'h0)] : ($unsigned((8'ha7)) ?
                      ($signed(reg419) ?
                          (forvar477 >>> reg448) : (~reg416)) : {(reg515 >>> reg483),
                          reg440})));
            end
          if ((reg397[(3'h4):(2'h3)] ?
              ($signed($unsigned({forvar407, reg498})) ?
                  $unsigned(reg482[(4'hb):(2'h2)]) : $signed(($signed(reg434) >> $unsigned(forvar449)))) : $unsigned(reg492)))
            begin
              reg518 = $unsigned($signed(((^~(reg487 ?
                  reg438 : reg420)) <= (!reg464[(3'h4):(1'h1)]))));
              reg519 <= $signed(({$unsigned((reg392 ? forvar407 : reg429)),
                      reg438} ?
                  ($unsigned(reg506[(4'hb):(1'h1)]) >> reg421) : $unsigned(reg426[(3'h5):(1'h1)])));
            end
          else
            begin
              reg518 <= (~&$signed($signed({$unsigned(reg438), (8'hbc)})));
              reg519 = ($signed(forvar512[(1'h0):(1'h0)]) ?
                  $signed($unsigned(reg435)) : (reg408[(3'h4):(1'h0)] ?
                      reg476[(1'h0):(1'h0)] : reg429[(1'h0):(1'h0)]));
              reg520 = (~reg448);
              reg521 <= ("Hp99yRzV" >> (($signed($unsigned(reg398)) && ($unsigned(reg408) ?
                  $unsigned(reg405) : {reg421})) + reg476[(4'ha):(4'h9)]));
            end
        end
      reg522 <= {reg496,
          ($signed((reg472 ?
                  $signed(reg491) : (reg423 ? forvar446 : (8'hb6)))) ?
              $unsigned(((|reg434) ?
                  {(8'h9e), (8'ha5)} : $signed(reg497))) : (-"6rr2ou9P"))};
    end
  always
    @(posedge clk) begin
      reg523 = $unsigned(reg422[(4'hc):(4'hb)]);
      if (((~^reg508) ?
          reg445 : (reg522 != ((|reg400) ?
              forvar477[(1'h0):(1'h0)] : $unsigned(((8'h9e) ?
                  reg461 : reg413))))))
        begin
          for (forvar524 = (1'h0); (forvar524 < (3'h4)); forvar524 = (forvar524 + (1'h1)))
            begin
              reg525 <= $signed($unsigned(reg510[(2'h2):(1'h1)]));
              reg526 = (({wire388[(4'h9):(4'h9)],
                      ((reg505 ^ reg465) ? reg428 : $signed((7'h42)))} ?
                  (~|$signed($signed(reg481))) : (~^forvar495[(2'h3):(1'h0)])) || (wire386 ?
                  (-($unsigned(forvar432) == $unsigned(forvar429))) : (~|{forvar493})));
              reg527 <= $unsigned({$signed(($unsigned(reg510) ?
                      $unsigned(reg429) : ((8'hbc) ? forvar471 : forvar514)))});
            end
          if (reg395)
            begin
              reg528 = "n0VFNvSfuRkiyivOxTMS";
              reg529 = $signed($unsigned(reg448));
            end
          else
            begin
              reg528 = reg465;
              reg529 = $signed(reg432[(2'h2):(2'h2)]);
              reg530 <= ($unsigned((forvar503 ?
                  $unsigned($unsigned(reg428)) : ((reg475 >> reg411) || (~reg420)))) ^~ $unsigned($signed($unsigned((forvar471 ?
                  (8'hbe) : forvar438)))));
              reg531 = reg456[(4'h8):(3'h7)];
            end
          if ((reg431[(1'h0):(1'h0)] <= reg413[(3'h5):(1'h1)]))
            begin
              reg532 <= $signed($signed($signed(forvar457)));
              reg533 <= $signed(($signed(($signed(reg441) ?
                      $signed(forvar432) : $signed((8'hbc)))) ?
                  $signed(reg405[(3'h6):(3'h6)]) : ((8'ha6) ?
                      reg394[(4'h8):(1'h0)] : (reg489[(2'h3):(2'h2)] ?
                          reg417[(3'h4):(2'h2)] : $unsigned((8'ha8))))));
              reg534 <= ($signed({reg429[(2'h2):(2'h2)],
                  ((!reg420) ?
                      (!(8'hbd)) : $signed(reg522))}) >= $signed((({wire386} & (^(8'hb1))) ?
                  {(8'hbd)} : $signed((reg479 | reg472)))));
              reg535 <= (~(reg408 ? forvar451 : (^reg434[(1'h1):(1'h0)])));
            end
          else
            begin
              reg532 <= $signed({(reg463[(4'hf):(4'h8)] ?
                      ((reg474 ? reg467 : reg434) & $signed(reg399)) : reg450),
                  (reg411 + $signed("hTPNRpkCI697eN"))});
              reg533 <= (reg494[(4'h8):(3'h7)] == $signed($unsigned((~|(reg415 ?
                  forvar511 : (8'ha8))))));
            end
        end
      else
        begin
          if ($unsigned(((~|($unsigned(reg397) && $unsigned(reg480))) | (~forvar460[(3'h5):(3'h5)]))))
            begin
              reg524 <= forvar495[(2'h3):(2'h3)];
              reg525 <= ((^(((-reg415) - (reg485 ? reg519 : reg445)) ?
                      ((reg401 >= reg442) ?
                          (^~(8'ha4)) : (reg421 ?
                              wire500 : (8'ha8))) : reg408)) ?
                  $signed((wire387[(4'hc):(1'h0)] ?
                      {(reg517 << forvar493)} : (^~{(8'h9c)}))) : (reg398[(2'h2):(2'h2)] ?
                      {$unsigned($unsigned(reg490))} : ($signed((reg517 ?
                          forvar393 : reg397)) ^~ reg402[(3'h6):(3'h6)])));
            end
          else
            begin
              reg524 = reg433[(1'h1):(1'h1)];
              reg525 = "sM84z9MwgUiAqt5";
              reg526 <= $unsigned($unsigned(reg419[(2'h3):(2'h2)]));
              reg527 <= (~|$unsigned(reg463));
              reg528 = (8'hb5);
            end
          for (forvar529 = (1'h0); (forvar529 < (3'h4)); forvar529 = (forvar529 + (1'h1)))
            begin
              reg530 <= $signed($unsigned((((8'hb4) ?
                  (forvar418 ?
                      forvar447 : reg399) : (reg496 ^~ (8'hbc))) == {(forvar438 ?
                      reg436 : reg458),
                  (~^reg524)})));
              reg531 <= (reg527 < reg430);
              reg532 <= ((($signed($unsigned(reg423)) ?
                  $unsigned((reg455 ?
                      forvar437 : reg452)) : $unsigned($unsigned(reg475))) <= ($signed(reg531) ?
                  forvar507 : (forvar418[(1'h0):(1'h0)] ?
                      forvar478[(2'h3):(2'h2)] : reg463[(4'h8):(3'h6)]))) - (reg428[(4'hc):(4'ha)] ?
                  reg397 : $signed({"GW", (forvar529 ? reg513 : reg435)})));
            end
          for (forvar533 = (1'h0); (forvar533 < (1'h1)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 = reg409;
            end
          reg535 = (8'hbf);
        end
      if (reg443)
        begin
          reg536 <= ((!reg438) <<< reg417);
        end
      else
        begin
          reg536 <= (((&forvar457[(4'ha):(3'h5)]) || ({(reg436 ?
                      (8'ha1) : forvar533),
                  {reg506, reg485}} ?
              $signed((reg409 >= (8'hae))) : reg461)) * $signed($signed((7'h44))));
          for (forvar537 = (1'h0); (forvar537 < (1'h1)); forvar537 = (forvar537 + (1'h1)))
            begin
              reg538 <= reg427[(1'h1):(1'h1)];
              reg539 <= wire499[(4'h9):(4'h9)];
              reg540 <= ({$signed(reg400),
                  {$signed($signed(reg517)),
                      reg529}} >> ((8'h9d) >> forvar477));
              reg541 = {$unsigned(reg439[(2'h2):(1'h0)])};
            end
          for (forvar542 = (1'h0); (forvar542 < (2'h2)); forvar542 = (forvar542 + (1'h1)))
            begin
              reg543 <= ($signed((~|$signed(reg529[(2'h2):(1'h0)]))) ?
                  ($signed((|reg450)) + $unsigned({forvar446,
                      "DUUvO11crwF6ag"})) : reg416[(1'h0):(1'h0)]);
              reg544 <= $unsigned({($unsigned(forvar502) ?
                      ((reg440 ? reg433 : (8'hae)) ?
                          (reg535 ?
                              reg445 : wire388) : reg430[(3'h5):(2'h3)]) : ((forvar412 * reg497) ?
                          reg455 : reg444)),
                  $unsigned((((8'haf) ?
                      reg432 : reg440) << (forvar503 >= forvar451)))});
              reg545 <= ((reg414 ?
                  ((|forvar457[(1'h1):(1'h1)]) != $signed(reg465)) : forvar446[(4'hc):(4'h8)]) && {({(~|wire388),
                          reg531[(4'ha):(1'h1)]} ?
                      ((forvar418 ?
                          (7'h44) : forvar542) <<< forvar441[(3'h6):(2'h3)]) : reg400[(5'h14):(4'hd)]),
                  forvar429});
              reg546 = ((($unsigned((reg505 == reg394)) ?
                      (8'hbd) : reg408[(2'h3):(1'h1)]) && (forvar542 & forvar478[(2'h3):(1'h1)])) ?
                  {(reg543 >= {forvar437[(4'ha):(4'h9)],
                          (wire389 ? forvar478 : (8'hae))}),
                      $unsigned((!(forvar495 ?
                          reg393 : reg424)))} : $signed((-((-forvar507) << $signed((8'hb7))))));
              reg547 = reg532[(2'h3):(2'h3)];
            end
          reg548 <= $unsigned(wire500[(2'h3):(2'h3)]);
          for (forvar549 = (1'h0); (forvar549 < (2'h3)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= {(&$unsigned(($signed((8'h9d)) >>> $signed((8'hb6))))),
                  $unsigned(forvar524[(1'h1):(1'h1)])};
              reg551 <= (wire388[(4'hc):(1'h1)] << ($signed(reg445[(3'h5):(1'h1)]) ?
                  reg529[(3'h5):(2'h2)] : (($unsigned(forvar514) >>> forvar537) ?
                      $signed((^forvar524)) : ($signed(reg489) - forvar502))));
              reg552 = reg454;
              reg553 = $unsigned(forvar429[(1'h0):(1'h0)]);
              reg554 <= $signed($unsigned($signed({$unsigned(reg419)})));
            end
        end
      reg555 <= {$unsigned({reg410})};
      reg556 <= (!($unsigned((~|reg547[(4'he):(4'hc)])) < (~^(forvar502[(5'h11):(3'h7)] * (&reg535)))));
    end
  always
    @(posedge clk) begin
      reg557 = ($signed(reg396) ?
          reg474 : (($unsigned({reg461}) ?
                  "NV" : (reg437[(5'h14):(4'hd)] ?
                      ((7'h44) == reg475) : reg526)) ?
              (((reg506 ? reg551 : reg438) <= $unsigned(forvar524)) ?
                  ({reg392, reg532} ^~ "d4bnP") : {(~(8'ha5)),
                      (!reg394)}) : $unsigned((forvar437 ?
                  {reg431, wire387} : (~|reg433)))));
      if ($unsigned(((($unsigned(reg463) == (-reg548)) ?
          reg557 : ("LnYuncUQCq5xPTBhLi" ?
              reg517[(4'hf):(4'hb)] : (wire390 < reg509))) < reg455)))
        begin
          for (forvar558 = (1'h0); (forvar558 < (2'h2)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 <= (8'ha0);
              reg560 = (reg522[(2'h2):(2'h2)] ? reg496 : reg551);
              reg561 <= $signed(({(~reg462),
                  $unsigned((reg528 > reg433))} != $signed((|(reg455 ?
                  forvar512 : wire501)))));
              reg562 <= (reg557[(2'h2):(1'h0)] >= ($unsigned(((forvar558 ^~ (8'hbe)) ?
                  $signed((8'hb5)) : (reg474 < reg559))) + reg396[(1'h0):(1'h0)]));
              reg563 <= reg545;
            end
          reg564 = $signed(((forvar406[(2'h3):(2'h2)] * ($unsigned(reg483) ?
                  (reg536 ? reg523 : reg548) : $signed(reg521))) ?
              reg455[(3'h4):(2'h3)] : forvar503));
          reg565 <= forvar507[(3'h6):(2'h2)];
        end
      else
        begin
          for (forvar558 = (1'h0); (forvar558 < (1'h1)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 <= (^~((reg485 != (reg479[(5'h11):(4'ha)] <= $signed((8'hbb)))) ?
                  {($unsigned((8'ha7)) ?
                          (|reg428) : (|forvar537))} : (((reg564 ?
                              reg508 : forvar471) ?
                          $signed((7'h41)) : reg508) ?
                      ((+forvar478) ?
                          (|reg556) : (reg539 ?
                              reg513 : reg474)) : reg476[(3'h7):(3'h7)])));
            end
          for (forvar560 = (1'h0); (forvar560 < (2'h3)); forvar560 = (forvar560 + (1'h1)))
            begin
              reg561 <= (|reg397[(2'h3):(1'h0)]);
              reg562 = reg524[(4'hc):(4'ha)];
              reg563 <= ($unsigned(reg561[(3'h6):(3'h5)]) <<< ((reg461 * (|$signed(reg544))) ?
                  $signed(forvar488[(3'h4):(1'h1)]) : forvar437));
              reg564 <= (~&$signed({(reg565[(3'h4):(3'h4)] ?
                      $signed(reg554) : forvar451[(3'h4):(1'h0)])}));
            end
        end
      for (forvar566 = (1'h0); (forvar566 < (1'h0)); forvar566 = (forvar566 + (1'h1)))
        begin
          for (forvar567 = (1'h0); (forvar567 < (2'h2)); forvar567 = (forvar567 + (1'h1)))
            begin
              reg568 <= {($signed($unsigned($unsigned(forvar566))) ?
                      (((forvar542 >>> forvar428) ?
                              $unsigned(reg510) : $unsigned(forvar457)) ?
                          reg496[(3'h4):(3'h4)] : reg401) : $unsigned($signed($unsigned(reg479))))};
              reg569 <= "066xSp36HM";
              reg570 <= (+$signed((~^(reg424 ?
                  reg440 : (reg483 ? reg552 : reg530)))));
              reg571 = ($signed(reg505[(2'h3):(2'h2)]) ?
                  (~&reg394) : (~^($unsigned((8'ha2)) ?
                      forvar451 : $signed(reg531))));
            end
          for (forvar572 = (1'h0); (forvar572 < (2'h2)); forvar572 = (forvar572 + (1'h1)))
            begin
              reg573 = {$signed($signed({(reg530 << forvar449)})),
                  {{forvar512,
                          ((forvar478 ? reg414 : reg545) ?
                              reg550[(4'hf):(2'h2)] : (^reg428))},
                      reg531[(4'hb):(4'ha)]}};
              reg574 <= wire500;
              reg575 <= $signed(reg419[(1'h0):(1'h0)]);
            end
          reg576 <= {forvar460[(3'h6):(1'h1)],
              (({$unsigned(reg414)} ?
                  reg401[(3'h5):(2'h3)] : (-(reg482 ?
                      forvar447 : reg487))) * reg463[(4'hb):(4'hb)])};
        end
    end
  assign wire577 = $unsigned((reg452 != (+{$signed(reg504),
                       $unsigned(reg468)})));
  assign wire578 = (-(~reg400[(5'h10):(3'h6)]));
  always
    @(posedge clk) begin
      for (forvar579 = (1'h0); (forvar579 < (2'h3)); forvar579 = (forvar579 + (1'h1)))
        begin
          if ({(&{((8'hb9) ? reg528[(4'h8):(2'h2)] : (forvar432 > reg453))})})
            begin
              reg580 <= ((reg482[(3'h6):(1'h0)] + reg392) ~^ $unsigned((($signed(reg554) > {reg485}) < $signed($signed((8'hb3))))));
              reg581 <= ($signed(reg489[(4'hc):(3'h5)]) < forvar495[(3'h6):(2'h3)]);
              reg582 <= reg490[(4'ha):(3'h6)];
              reg583 = ((($signed((forvar457 >>> reg563)) ~^ (+((8'hab) >> (8'ha3)))) ?
                      $signed(((~|reg575) >> reg557)) : $unsigned((reg481[(3'h4):(2'h2)] ?
                          reg473[(2'h3):(1'h0)] : forvar451))) ?
                  reg458[(1'h0):(1'h0)] : $signed({$unsigned((~|forvar429))}));
              reg584 = ($signed(((^((8'ha3) + forvar566)) | forvar542)) ?
                  wire578 : (((8'hbf) >= reg546[(5'h10):(4'h9)]) <= reg394[(4'ha):(1'h0)]));
            end
          else
            begin
              reg580 <= $signed($signed(($signed($unsigned(reg494)) << "JIEdLL5YgGGL8Pi0zS6e")));
              reg581 <= (|reg522);
            end
          reg585 <= $unsigned(reg551);
          reg586 = $signed($signed((reg576[(1'h0):(1'h0)] ?
              wire388[(5'h14):(4'hc)] : {{forvar466, (7'h44)},
                  $signed(reg520)})));
          for (forvar587 = (1'h0); (forvar587 < (1'h0)); forvar587 = (forvar587 + (1'h1)))
            begin
              reg588 <= {reg491[(1'h0):(1'h0)]};
              reg589 = $signed((^~(^{(reg494 ? reg454 : reg429)})));
              reg590 <= $signed(reg534);
              reg591 = "lfb5k8I8U";
              reg592 <= {(~^($signed(((8'ha9) ? reg486 : wire577)) ?
                      reg417 : reg531))};
            end
          for (forvar593 = (1'h0); (forvar593 < (1'h1)); forvar593 = (forvar593 + (1'h1)))
            begin
              reg594 = ($signed((^reg456)) <<< "aD");
              reg595 <= (-$unsigned((^~$unsigned({forvar529}))));
              reg596 <= $unsigned(reg448);
              reg597 <= $unsigned(((^~forvar447) ?
                  (~^(reg420 ?
                      (reg496 ?
                          wire577 : reg522) : (reg430 + reg396))) : (&(forvar507[(5'h10):(5'h10)] ?
                      (reg459 ? reg509 : reg521) : ((7'h41) ?
                          reg430 : (8'h9e))))));
            end
        end
      reg598 <= ((reg416[(3'h5):(3'h4)] ?
              reg519 : (reg582[(4'ha):(4'h8)] + $unsigned($unsigned(reg592)))) ?
          reg474[(3'h4):(1'h0)] : reg492);
      reg599 = reg556[(3'h5):(1'h0)];
      for (forvar600 = (1'h0); (forvar600 < (1'h0)); forvar600 = (forvar600 + (1'h1)))
        begin
          reg601 <= (&((~&$signed($unsigned(reg439))) << reg551[(1'h0):(1'h0)]));
          reg602 <= (8'ha1);
          reg603 = $unsigned(((reg594[(3'h5):(1'h1)] - ($signed(reg394) < {(8'haf)})) - (~&(~|forvar587[(4'h9):(3'h4)]))));
          for (forvar604 = (1'h0); (forvar604 < (2'h3)); forvar604 = (forvar604 + (1'h1)))
            begin
              reg605 <= $unsigned((8'hb3));
              reg606 <= {((forvar511[(3'h5):(2'h2)] ^~ reg445[(4'hb):(1'h0)]) ?
                      reg405[(4'h8):(3'h6)] : (((reg433 ?
                              (8'hae) : forvar495) & {reg533, (8'hb2)}) ?
                          ({reg505} >>> reg397[(2'h2):(1'h1)]) : "xLOQT6m0TaL7izPCuE9K"))};
              reg607 = reg479[(4'hc):(1'h0)];
            end
        end
      if (((&$unsigned(reg505[(1'h1):(1'h1)])) ?
          ($unsigned({$unsigned(reg394)}) > $signed((~|(^(8'ha5))))) : $unsigned((|reg392))))
        begin
          reg608 = (wire389 ^~ reg596);
          for (forvar609 = (1'h0); (forvar609 < (2'h2)); forvar609 = (forvar609 + (1'h1)))
            begin
              reg610 <= $unsigned(reg551);
              reg611 <= ((+$signed((!(~&forvar609)))) ?
                  ({$unsigned((reg445 ? reg556 : reg426)), forvar447} ?
                      {{{forvar433},
                              (reg465 ?
                                  forvar609 : reg515)}} : $unsigned(reg561)) : ($unsigned(reg585[(3'h5):(2'h3)]) >= {reg413[(3'h5):(3'h4)]}));
            end
        end
      else
        begin
          reg608 <= reg437;
          for (forvar609 = (1'h0); (forvar609 < (2'h2)); forvar609 = (forvar609 + (1'h1)))
            begin
              reg610 <= ((reg571[(3'h6):(1'h1)] - $unsigned(reg601[(1'h1):(1'h0)])) ?
                  (+(reg491[(3'h4):(2'h2)] | (reg413 == (~|(8'h9e))))) : reg551);
              reg611 = {(~&(reg486[(3'h5):(2'h3)] ?
                      (!{reg590, reg476}) : ((reg563 ? reg527 : (8'ha0)) ?
                          (wire388 * reg458) : {reg498})))};
              reg612 <= "RKlx4bY2ng6JN2G";
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar613 = (1'h0); (forvar613 < (1'h0)); forvar613 = (forvar613 + (1'h1)))
        begin
          for (forvar614 = (1'h0); (forvar614 < (3'h4)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 <= reg535;
              reg616 <= "2eQ5w21GOBr5huXIx";
              reg617 <= forvar457;
              reg618 = reg539;
              reg619 = {forvar604[(4'ha):(3'h7)]};
            end
        end
      reg620 <= $signed(forvar537);
    end
  assign wire621 = (!$unsigned(reg564[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      for (forvar622 = (1'h0); (forvar622 < (2'h2)); forvar622 = (forvar622 + (1'h1)))
        begin
          reg623 <= ((reg430[(3'h6):(2'h2)] + (~(8'hb1))) ?
              reg557[(1'h1):(1'h1)] : $signed((-reg591)));
          reg624 = reg562;
          reg625 <= $signed((reg610[(4'he):(2'h2)] == (reg535[(4'ha):(2'h3)] >> (~{(8'hbd),
              (8'hb8)}))));
        end
      if ((wire386 ? $unsigned($signed($signed(forvar406))) : (~^forvar437)))
        begin
          reg626 = (reg580[(5'h14):(3'h4)] && ($signed(($unsigned(reg573) ?
                  {reg548} : $unsigned(forvar478))) ?
              reg409 : $signed(forvar600)));
          reg627 <= "ZNV93R";
          for (forvar628 = (1'h0); (forvar628 < (1'h1)); forvar628 = (forvar628 + (1'h1)))
            begin
              reg629 <= $signed($unsigned(reg589[(2'h2):(1'h0)]));
            end
          for (forvar630 = (1'h0); (forvar630 < (1'h0)); forvar630 = (forvar630 + (1'h1)))
            begin
              reg631 <= {"Z8SM1l9293XQk0TcfZPa"};
            end
          reg632 <= reg522[(1'h1):(1'h0)];
        end
      else
        begin
          reg626 <= $signed($signed({(((8'had) ? (8'had) : reg564) & reg416)}));
        end
      if ("pZ1YpbEbQA7d5Bil")
        begin
          reg633 <= reg557;
          for (forvar634 = (1'h0); (forvar634 < (2'h2)); forvar634 = (forvar634 + (1'h1)))
            begin
              reg635 = (reg485[(3'h4):(1'h1)] && {reg491[(2'h3):(1'h0)],
                  "1hp1g8JfAZXi902Ef"});
              reg636 = $unsigned($unsigned(((~^forvar542[(1'h1):(1'h1)]) ?
                  $signed((|reg599)) : (~&{reg420}))));
              reg637 = reg490[(3'h4):(1'h0)];
              reg638 <= (reg532[(2'h3):(2'h3)] ?
                  (~(((reg632 >= reg424) ?
                      reg632[(3'h7):(3'h5)] : $unsigned(wire500)) - reg538)) : $signed((((reg625 && reg560) ?
                      (reg423 - reg421) : (reg625 - (8'hac))) ^~ {$unsigned(reg633)})));
              reg639 = (8'ha2);
            end
          reg640 = {$unsigned("kMQ"), {(!$unsigned({forvar604}))}};
        end
      else
        begin
          reg633 = reg439;
        end
      for (forvar641 = (1'h0); (forvar641 < (2'h3)); forvar641 = (forvar641 + (1'h1)))
        begin
          reg642 <= $signed($unsigned($signed(forvar512)));
          reg643 = ($signed($signed(forvar558)) <= $unsigned(reg448));
          if ((8'ha0))
            begin
              reg644 <= $signed(wire387);
              reg645 = reg396;
              reg646 <= reg504;
              reg647 <= (($signed($signed((!forvar587))) ?
                  $signed(($unsigned(reg588) | (reg397 < forvar628))) : reg433[(1'h0):(1'h0)]) << $unsigned($signed(($signed(forvar542) ?
                  (8'hbd) : {(8'hae), forvar447}))));
              reg648 <= forvar542;
            end
          else
            begin
              reg644 <= ((+(-$signed({reg405,
                  forvar533}))) <= $unsigned($signed("dKoUfB")));
              reg645 = (forvar634[(2'h2):(1'h1)] ?
                  (((8'had) + {(reg576 | reg631)}) ?
                      (reg461[(4'hb):(2'h3)] ?
                          (8'hbb) : (~&{reg399,
                              (8'hbe)})) : reg648[(1'h1):(1'h0)]) : {$unsigned($signed((reg439 ?
                          (8'hbc) : reg560))),
                      (-$unsigned(reg569))});
              reg646 = $signed(reg482[(4'hc):(1'h0)]);
              reg647 <= ($signed((forvar393[(1'h0):(1'h0)] ?
                      (reg508[(3'h5):(1'h0)] ?
                          $signed(wire578) : (+reg408)) : forvar429)) ?
                  ($unsigned((|(reg594 > forvar477))) ?
                      {(^$unsigned(reg394)),
                          $unsigned("omH30eSbrm")} : $unsigned(reg574[(3'h5):(1'h0)])) : (^~$unsigned($unsigned($signed(reg510)))));
              reg648 <= (&($signed($signed({reg505})) ?
                  $signed(forvar433) : ($signed("BmOFL") & ($unsigned(reg602) == (reg561 ?
                      (8'ha5) : reg598)))));
            end
          if ("08Mhh8AYz")
            begin
              reg649 = {((+$unsigned($signed(reg633))) ?
                      $unsigned(reg574) : {(reg626 & (^~forvar466)),
                          ((^~(8'ha8)) <= {(8'h9e), wire621})}),
                  reg494[(2'h3):(1'h1)]};
              reg650 <= $unsigned((^($signed({reg440,
                  reg647}) >>> reg485[(4'h8):(1'h1)])));
              reg651 <= $unsigned($unsigned($signed((+"TEXDV1e49vVAwgkrbG0"))));
            end
          else
            begin
              reg649 <= (^$unsigned((8'hb6)));
              reg650 <= $unsigned($signed($signed(forvar471[(1'h1):(1'h0)])));
              reg651 <= ((!reg445) ?
                  {(($unsigned(reg525) && reg498) ?
                          (8'hb7) : ("plrDlIxzBt4IY" | reg524[(5'h12):(3'h6)]))} : (+reg618));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar652 = (1'h0); (forvar652 < (2'h2)); forvar652 = (forvar652 + (1'h1)))
        begin
          for (forvar653 = (1'h0); (forvar653 < (3'h4)); forvar653 = (forvar653 + (1'h1)))
            begin
              reg654 <= forvar511[(2'h2):(1'h0)];
              reg655 = $unsigned(forvar524[(1'h0):(1'h0)]);
              reg656 <= ((reg588 ? "ViLGKFFnrp4" : reg643[(2'h2):(1'h1)]) ?
                  $unsigned(forvar393) : $signed({$signed(reg642[(4'h9):(3'h4)])}));
              reg657 <= "S";
            end
          for (forvar658 = (1'h0); (forvar658 < (3'h4)); forvar658 = (forvar658 + (1'h1)))
            begin
              reg659 = (reg497 <<< {($signed((&reg469)) ?
                      {(reg603 ? reg556 : reg393)} : wire389[(5'h14):(4'hd)]),
                  forvar393});
              reg660 <= (-((reg523 ?
                      (reg581 >>> (~&reg404)) : ($signed(reg455) | (reg554 ?
                          reg416 : forvar451))) ?
                  ($signed((-forvar641)) ?
                      ($signed(reg465) ?
                          forvar630[(2'h2):(1'h0)] : reg456) : reg414) : ($signed((+forvar429)) ?
                      $unsigned(reg601[(1'h0):(1'h0)]) : (((8'ha5) << forvar572) - forvar451))));
            end
          reg661 <= reg504;
          if ((!(8'h9e)))
            begin
              reg662 <= {"ImZO"};
              reg663 = (+(|(~&"G6fhNaD3qEUZe7")));
              reg664 <= ($unsigned($unsigned(((~forvar406) ?
                  {(8'hb5)} : reg536[(3'h7):(3'h7)]))) == forvar567[(4'h9):(4'h8)]);
            end
          else
            begin
              reg662 = $signed($signed(($unsigned(reg430) ?
                  (~|$unsigned(reg539)) : reg413[(4'he):(4'h8)])));
              reg663 <= "hnq1Pp";
              reg664 = $signed($unsigned($signed(reg454)));
              reg665 <= reg560[(4'hf):(2'h3)];
            end
          for (forvar666 = (1'h0); (forvar666 < (2'h3)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 <= reg602[(4'hb):(3'h5)];
              reg668 = $signed($signed((!{(reg421 ? reg586 : forvar593)})));
              reg669 <= $signed($unsigned(reg586[(3'h4):(2'h2)]));
              reg670 <= $unsigned((reg434[(4'hb):(3'h7)] ?
                  reg392[(3'h4):(1'h1)] : ($unsigned((!(7'h40))) ?
                      (((8'haf) ^~ forvar502) ~^ {reg571}) : $signed({reg565,
                          forvar653}))));
            end
        end
      reg671 = {forvar488[(1'h0):(1'h0)]};
      reg672 <= ($unsigned(({(|forvar502),
          $signed(forvar567)} < reg650[(1'h0):(1'h0)])) | ((+"9bco3GE") ?
          $unsigned($signed(reg522)) : {reg627[(2'h2):(1'h1)],
              ($unsigned((8'hb4)) ? (7'h41) : ((8'ha9) - reg396))}));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module326
#( parameter param381 = (^~(~^(&((!(8'ha2)) && (+(8'ha8))))))
, parameter param382 = ((((!param381) ? (^~(~&param381)) : param381) & (&(param381 >>> (param381 ? param381 : param381)))) ? (&(((param381 != param381) ? ((8'haf) > param381) : (param381 - param381)) ? (((8'hb3) ^~ param381) ? param381 : (!param381)) : ({param381} ? param381 : param381))) : ((+(~&(|param381))) ? {(param381 ? (~&param381) : param381)} : (-(((8'h9c) ? param381 : param381) ^ param381)))) )
(y, clk, wire331, wire330, wire329, wire328, wire327);
  output wire [(32'h268):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire331;
  input wire signed [(3'h5):(1'h0)] wire330;
  input wire signed [(3'h7):(1'h0)] wire329;
  input wire signed [(4'h8):(1'h0)] wire328;
  input wire [(3'h5):(1'h0)] wire327;
  wire [(4'hb):(1'h0)] wire380;
  reg [(5'h11):(1'h0)] reg379 = (1'h0);
  reg [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar377 = (1'h0);
  reg [(3'h4):(1'h0)] reg376 = (1'h0);
  wire [(3'h5):(1'h0)] wire375;
  reg signed [(4'hf):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg373 = (1'h0);
  reg [(5'h10):(1'h0)] reg372 = (1'h0);
  reg [(4'hd):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg369 = (1'h0);
  reg [(5'h15):(1'h0)] forvar368 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg367 = (1'h0);
  reg [(4'ha):(1'h0)] reg366 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg365 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg364 = (1'h0);
  reg [(4'hf):(1'h0)] reg363 = (1'h0);
  reg [(4'hb):(1'h0)] forvar362 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg361 = (1'h0);
  reg [(4'hd):(1'h0)] reg360 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg359 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg358 = (1'h0);
  reg [(5'h11):(1'h0)] reg357 = (1'h0);
  reg [(4'hd):(1'h0)] forvar356 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg355 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire354;
  wire [(5'h14):(1'h0)] wire353;
  wire signed [(4'he):(1'h0)] wire352;
  wire [(4'hc):(1'h0)] wire351;
  wire signed [(4'hd):(1'h0)] wire350;
  wire [(3'h7):(1'h0)] wire349;
  reg [(4'he):(1'h0)] reg348 = (1'h0);
  reg [(5'h12):(1'h0)] reg347 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg346 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] reg344 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar343 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg341 = (1'h0);
  reg [(3'h4):(1'h0)] forvar340 = (1'h0);
  reg [(5'h15):(1'h0)] reg339 = (1'h0);
  reg [(5'h13):(1'h0)] forvar338 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar339 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg337 = (1'h0);
  reg [(4'hb):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg334 = (1'h0);
  reg [(3'h7):(1'h0)] reg333 = (1'h0);
  reg [(5'h15):(1'h0)] forvar332 = (1'h0);
  assign y = {wire380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 wire375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 forvar368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 forvar356,
                 reg355,
                 wire354,
                 wire353,
                 wire352,
                 wire351,
                 wire350,
                 wire349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 forvar343,
                 reg342,
                 reg341,
                 forvar340,
                 reg339,
                 forvar338,
                 reg340,
                 forvar339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 forvar332,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned(((wire330 ?
          $unsigned($unsigned((8'haa))) : wire331) < (wire331 ?
          ($signed(wire331) ~^ (wire328 == wire327)) : ((~wire328) ?
              ((8'hb1) ? wire330 : wire327) : wire331[(2'h3):(2'h2)])))))
        begin
          for (forvar332 = (1'h0); (forvar332 < (1'h1)); forvar332 = (forvar332 + (1'h1)))
            begin
              reg333 <= (wire330[(2'h2):(2'h2)] << (8'hba));
              reg334 = $signed(wire331[(4'h9):(2'h2)]);
              reg335 <= {"Qaxb5e", reg334[(2'h3):(1'h0)]};
              reg336 <= wire330[(3'h5):(1'h0)];
            end
          if (reg334[(4'hb):(1'h0)])
            begin
              reg337 <= $signed((!(((-wire327) * (8'ha1)) | $unsigned((wire328 > (8'had))))));
            end
          else
            begin
              reg337 = ((reg335 || (~$signed($unsigned(wire327)))) ?
                  $signed(((((8'hbb) ?
                      (7'h43) : reg336) | wire331[(4'hb):(1'h0)]) ^~ (^$signed(wire330)))) : (($unsigned($signed(wire331)) ?
                          ($unsigned(wire331) ? (8'hb5) : wire327) : wire329) ?
                      $signed((~reg335[(3'h5):(2'h2)])) : wire328[(2'h3):(2'h2)]));
              reg338 = (wire328 ?
                  reg334[(1'h1):(1'h0)] : $signed(($signed((8'ha5)) > wire329)));
            end
          for (forvar339 = (1'h0); (forvar339 < (1'h0)); forvar339 = (forvar339 + (1'h1)))
            begin
              reg340 = $unsigned((~&(reg335 ?
                  wire331 : (wire331[(2'h3):(1'h1)] < wire327))));
            end
        end
      else
        begin
          for (forvar332 = (1'h0); (forvar332 < (3'h4)); forvar332 = (forvar332 + (1'h1)))
            begin
              reg333 = (8'hbe);
              reg334 <= $signed($signed(reg333[(1'h1):(1'h1)]));
              reg335 = wire328;
              reg336 = $signed(({((&(8'hb1)) <<< (^~reg335))} ?
                  {((wire330 ? (8'hbb) : reg340) + wire330),
                      forvar332} : $unsigned($signed($unsigned(reg335)))));
              reg337 = ((+$unsigned($signed((reg337 ?
                  wire331 : reg333)))) <<< $signed($unsigned((!(forvar339 ?
                  reg337 : (8'hbf))))));
            end
          for (forvar338 = (1'h0); (forvar338 < (2'h2)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 <= (^~$unsigned({($signed((7'h40)) ? (^~reg334) : wire328),
                  $signed((-forvar339))}));
            end
          for (forvar340 = (1'h0); (forvar340 < (2'h2)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 = "9ef1kb5HEt";
              reg342 <= reg335[(4'ha):(3'h5)];
            end
          for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 = (~(~^reg335));
              reg345 <= forvar332[(5'h12):(4'hf)];
              reg346 = wire329;
              reg347 = {$signed($signed($signed(((7'h41) & wire330))))};
              reg348 = $signed($signed($unsigned($unsigned($signed(reg342)))));
            end
        end
    end
  assign wire349 = reg346;
  assign wire350 = ((8'hbd) ^~ wire329[(3'h4):(1'h1)]);
  assign wire351 = wire349;
  assign wire352 = (~^((^wire331[(4'ha):(2'h3)]) ?
                       (reg336[(2'h3):(2'h2)] ?
                           {reg345[(2'h2):(1'h1)],
                               $signed(reg348)} : (8'hb4)) : (reg337[(4'h9):(1'h1)] < {(wire327 ~^ reg348)})));
  assign wire353 = ((($signed((wire349 | wire327)) ?
                       $signed(wire328) : $unsigned(forvar338[(5'h11):(3'h5)])) && $signed(((wire351 & reg348) ?
                       reg333 : reg340[(1'h1):(1'h1)]))) > ((8'ha7) ?
                       (^(+(wire350 >>> reg333))) : forvar332[(5'h15):(4'h9)]));
  assign wire354 = (~|($unsigned((~|$signed(reg338))) ?
                       reg348 : $unsigned($signed(wire352))));
  always
    @(posedge clk) begin
      reg355 <= ((8'hb9) ?
          (!$unsigned("WykoHhSnfdcpu")) : $signed($signed(reg341[(5'h11):(1'h0)])));
      for (forvar356 = (1'h0); (forvar356 < (1'h0)); forvar356 = (forvar356 + (1'h1)))
        begin
          if (reg336[(3'h5):(3'h4)])
            begin
              reg357 = $unsigned(reg334[(5'h11):(5'h10)]);
            end
          else
            begin
              reg357 = ($unsigned((($signed(wire329) ?
                      (reg334 ~^ wire328) : $unsigned((7'h41))) ?
                  (((7'h43) >> reg339) ?
                      reg341 : (forvar339 ?
                          reg355 : forvar338)) : wire327)) ^~ (reg337[(2'h3):(2'h2)] ?
                  reg335 : (|(-(7'h40)))));
              reg358 = (8'hb5);
              reg359 = ("R98hpN7LXl4" ?
                  reg357 : (((reg344[(1'h0):(1'h0)] ^ wire329) ^~ (wire351[(1'h1):(1'h0)] & (~&reg340))) ?
                      reg342 : (!(8'hb3))));
              reg360 <= {{(((reg338 || (8'hba)) <<< (reg341 ?
                          reg345 : reg336)) ^~ $unsigned({forvar338, wire351})),
                      $unsigned(("YLCWH3f7EeEy7q" | ((8'h9f) ?
                          reg341 : reg333)))}};
              reg361 = ($unsigned($unsigned($signed((wire351 ?
                  reg358 : (8'hbd))))) <= reg333[(3'h4):(2'h3)]);
            end
          for (forvar362 = (1'h0); (forvar362 < (3'h4)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 = ((~|reg359) ?
                  (8'ha3) : $signed(((^~(reg355 + reg340)) ?
                      (&(+(8'hb5))) : wire350)));
              reg364 <= ($unsigned((((~|reg338) ?
                          $unsigned(reg358) : (+forvar339)) ?
                      reg334 : wire349[(3'h4):(2'h3)])) ?
                  reg336 : {($signed((reg347 ^ reg347)) ?
                          (+$signed(reg335)) : wire328[(1'h0):(1'h0)]),
                      $signed(((forvar340 ?
                          (8'hbb) : reg335) >= "iAaTHev9FwZsrqwIcJK"))});
              reg365 <= ((|(~wire327[(1'h0):(1'h0)])) - ((7'h42) ^~ (~|reg333[(3'h4):(1'h1)])));
              reg366 <= reg347;
              reg367 <= ($unsigned(reg363[(1'h0):(1'h0)]) ?
                  reg338[(2'h2):(1'h1)] : reg366[(3'h5):(2'h3)]);
            end
          for (forvar368 = (1'h0); (forvar368 < (2'h2)); forvar368 = (forvar368 + (1'h1)))
            begin
              reg369 = (-$signed(reg345));
              reg370 <= $signed($signed(reg333[(1'h0):(1'h0)]));
              reg371 <= $unsigned(({reg360} ?
                  $signed({(^wire354)}) : (reg338 ?
                      reg358[(1'h0):(1'h0)] : $signed($unsigned(wire351)))));
              reg372 <= (8'hb8);
              reg373 = (^(~|$signed((-(8'ha6)))));
            end
        end
      reg374 <= ((~&$signed($unsigned(reg358[(2'h2):(1'h0)]))) ?
          ((-((reg345 ? reg363 : (8'ha3)) ?
                  (reg369 == reg359) : (reg363 > wire328))) ?
              (((forvar362 ? (8'ha4) : reg355) ?
                      ((8'hb6) <<< reg347) : $signed(reg373)) ?
                  ({wire327} ?
                      reg366 : reg337) : $signed((-(8'hb5)))) : ((^(~^reg348)) ?
                  $signed(reg338) : (~|reg357))) : (~^$unsigned(((forvar343 ?
                  reg334 : reg345) ?
              (~forvar362) : $signed(reg369)))));
    end
  assign wire375 = reg337[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg376 <= "Eyo3SuDB";
      for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
        begin
          reg378 <= wire331[(1'h1):(1'h0)];
          reg379 <= $unsigned($signed($signed(reg366[(3'h6):(3'h6)])));
        end
    end
  assign wire380 = "BCU2tUEcMa";
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module204
#( parameter param319 = (~((~(&((7'h40) ? (7'h43) : (7'h43)))) || ((((8'ha7) >>> (8'haf)) && (~^(8'hae))) ? (((8'ha2) || (7'h40)) ? (^~(8'ha3)) : ((7'h44) ? (8'hb1) : (8'ha6))) : (((7'h42) ? (8'ha3) : (8'hb9)) | (!(8'ha2)))))) )
(y, clk, wire208, wire207, wire206, wire205);
  output wire [(32'h536):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire208;
  input wire signed [(4'h9):(1'h0)] wire207;
  input wire [(2'h2):(1'h0)] wire206;
  input wire [(5'h14):(1'h0)] wire205;
  reg [(3'h7):(1'h0)] reg318 = (1'h0);
  reg [(2'h3):(1'h0)] reg317 = (1'h0);
  reg [(2'h3):(1'h0)] forvar316 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg315 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg314 = (1'h0);
  reg [(4'hd):(1'h0)] reg313 = (1'h0);
  reg [(4'h9):(1'h0)] reg312 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar311 = (1'h0);
  reg [(4'hb):(1'h0)] reg310 = (1'h0);
  reg [(2'h3):(1'h0)] forvar305 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg309 = (1'h0);
  reg [(5'h13):(1'h0)] reg308 = (1'h0);
  reg [(5'h12):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg306 = (1'h0);
  reg [(2'h2):(1'h0)] reg305 = (1'h0);
  reg [(4'h9):(1'h0)] reg304 = (1'h0);
  reg [(4'hd):(1'h0)] reg303 = (1'h0);
  reg [(4'h9):(1'h0)] reg302 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg301 = (1'h0);
  reg [(4'he):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg299 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg297 = (1'h0);
  reg [(4'hd):(1'h0)] reg296 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg295 = (1'h0);
  reg [(4'he):(1'h0)] reg294 = (1'h0);
  reg [(3'h7):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar291 = (1'h0);
  reg [(4'ha):(1'h0)] reg290 = (1'h0);
  wire [(3'h6):(1'h0)] wire289;
  wire [(4'hb):(1'h0)] wire288;
  wire signed [(4'h9):(1'h0)] wire287;
  wire signed [(5'h15):(1'h0)] wire286;
  wire signed [(5'h10):(1'h0)] wire285;
  reg signed [(3'h4):(1'h0)] reg284 = (1'h0);
  reg [(5'h14):(1'h0)] reg283 = (1'h0);
  reg [(5'h14):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg281 = (1'h0);
  reg [(2'h3):(1'h0)] reg280 = (1'h0);
  reg [(5'h15):(1'h0)] forvar279 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar277 = (1'h0);
  reg [(4'hc):(1'h0)] reg276 = (1'h0);
  reg [(2'h3):(1'h0)] reg275 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg274 = (1'h0);
  reg [(5'h12):(1'h0)] reg273 = (1'h0);
  reg [(5'h12):(1'h0)] forvar272 = (1'h0);
  reg [(4'hd):(1'h0)] reg271 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar269 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg267 = (1'h0);
  reg [(4'ha):(1'h0)] forvar266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg265 = (1'h0);
  reg [(5'h15):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg263 = (1'h0);
  reg [(4'he):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg261 = (1'h0);
  reg [(3'h7):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg259 = (1'h0);
  reg [(4'h8):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar256 = (1'h0);
  reg [(4'hc):(1'h0)] forvar255 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire254;
  wire signed [(5'h15):(1'h0)] wire253;
  wire [(4'hb):(1'h0)] wire252;
  wire signed [(4'ha):(1'h0)] wire251;
  reg signed [(4'ha):(1'h0)] reg250 = (1'h0);
  reg [(3'h5):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg248 = (1'h0);
  reg [(2'h3):(1'h0)] reg247 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg245 = (1'h0);
  reg [(3'h4):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg243 = (1'h0);
  reg [(4'hf):(1'h0)] reg242 = (1'h0);
  reg signed [(4'he):(1'h0)] reg241 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg239 = (1'h0);
  reg [(4'hf):(1'h0)] forvar238 = (1'h0);
  reg [(4'ha):(1'h0)] forvar237 = (1'h0);
  reg [(4'hc):(1'h0)] reg236 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg234 = (1'h0);
  reg [(3'h7):(1'h0)] forvar233 = (1'h0);
  reg [(5'h10):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] reg228 = (1'h0);
  reg [(5'h10):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar223 = (1'h0);
  reg [(5'h14):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg219 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg218 = (1'h0);
  wire [(4'h8):(1'h0)] wire217;
  wire signed [(3'h4):(1'h0)] wire216;
  reg [(5'h10):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar214 = (1'h0);
  reg [(5'h14):(1'h0)] reg213 = (1'h0);
  reg signed [(4'he):(1'h0)] reg212 = (1'h0);
  reg [(4'he):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar210 = (1'h0);
  reg [(5'h13):(1'h0)] forvar209 = (1'h0);
  assign y = {reg318,
                 reg317,
                 forvar316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 forvar311,
                 reg310,
                 forvar305,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 forvar291,
                 reg290,
                 wire289,
                 wire288,
                 wire287,
                 wire286,
                 wire285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 forvar279,
                 reg278,
                 forvar277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 reg271,
                 reg270,
                 forvar269,
                 reg268,
                 reg267,
                 forvar266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 forvar256,
                 forvar255,
                 wire254,
                 wire253,
                 wire252,
                 wire251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 forvar238,
                 forvar237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 forvar223,
                 reg222,
                 reg221,
                 forvar220,
                 reg219,
                 reg218,
                 wire217,
                 wire216,
                 reg215,
                 forvar214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 forvar209,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar209 = (1'h0); (forvar209 < (1'h0)); forvar209 = (forvar209 + (1'h1)))
        begin
          for (forvar210 = (1'h0); (forvar210 < (1'h1)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= (wire208[(3'h7):(2'h2)] ?
                  (8'h9d) : $unsigned(($signed($unsigned(wire206)) <= ((wire206 != forvar209) ?
                      (wire208 ? forvar210 : wire206) : {forvar210}))));
              reg212 = $unsigned((((~|$signed(wire206)) ?
                      {$signed(forvar210)} : wire208) ?
                  (wire205 ? (8'hbd) : wire206) : reg211[(3'h7):(1'h0)]));
              reg213 <= forvar210[(2'h3):(2'h3)];
            end
          for (forvar214 = (1'h0); (forvar214 < (3'h4)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 = wire205[(5'h11):(3'h4)];
            end
        end
    end
  assign wire216 = reg211;
  assign wire217 = ((reg213 && reg213) ?
                       ($unsigned(((forvar210 ^~ wire205) >>> (wire205 ?
                           reg212 : forvar214))) ^ ({$signed(reg215)} > reg211)) : (8'hbf));
  always
    @(posedge clk) begin
      reg218 = (wire205[(4'hd):(1'h1)] ? forvar214 : wire208[(2'h2):(1'h0)]);
      reg219 = $unsigned((reg211[(1'h0):(1'h0)] ^ wire208[(3'h6):(1'h1)]));
      for (forvar220 = (1'h0); (forvar220 < (3'h4)); forvar220 = (forvar220 + (1'h1)))
        begin
          reg221 = wire205;
          reg222 <= wire208;
        end
      for (forvar223 = (1'h0); (forvar223 < (1'h1)); forvar223 = (forvar223 + (1'h1)))
        begin
          reg224 <= $signed(($unsigned(($signed(forvar209) ^~ {reg219,
                  wire205})) ?
              $unsigned(wire205) : (reg213 ?
                  ({(8'hb5), forvar220} >= reg212) : $unsigned((-wire205)))));
          if ($unsigned(reg213[(5'h11):(2'h2)]))
            begin
              reg225 = ((8'ha1) << (^~$unsigned({(~forvar214)})));
              reg226 = forvar214[(2'h3):(2'h2)];
              reg227 = reg221[(4'h9):(3'h4)];
              reg228 = ((~^(8'ha2)) ? wire217[(3'h4):(2'h3)] : wire207);
            end
          else
            begin
              reg225 = (+(($unsigned((|(8'ha7))) | reg219[(2'h2):(1'h0)]) - $unsigned((reg222[(4'ha):(4'h8)] ?
                  {forvar209} : (~^wire217)))));
            end
          reg229 <= (forvar210 ?
              $signed((^~("UFe10kK" ?
                  {forvar209,
                      forvar210} : wire207))) : $unsigned(((~|$unsigned(wire217)) == $unsigned($unsigned(reg213)))));
          reg230 <= (reg222 <= (reg225[(4'hf):(3'h4)] != $unsigned((~^{(8'hb3)}))));
        end
      if ((-($signed(forvar223) - (^~$unsigned((wire217 <= wire205))))))
        begin
          reg231 <= $signed(reg226);
        end
      else
        begin
          reg231 <= $unsigned(reg227[(3'h7):(2'h2)]);
          reg232 <= ($signed($signed(reg228[(2'h2):(1'h1)])) > ($signed($unsigned($signed((8'ha0)))) * $signed({$signed(reg231)})));
          for (forvar233 = (1'h0); (forvar233 < (2'h2)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 <= (forvar233[(3'h6):(1'h1)] <= ($unsigned("o") >>> reg213[(4'hd):(3'h6)]));
            end
          reg235 <= ((~forvar233) ?
              ((wire207 || $unsigned((!reg212))) ?
                  $signed((&forvar209[(4'hc):(2'h2)])) : reg222) : {(~&wire205),
                  (^reg232[(4'hf):(1'h1)])});
        end
    end
  always
    @(posedge clk) begin
      reg236 <= (+((wire206 ?
          $unsigned(reg226) : ($signed(reg235) != {forvar220})) > $signed(({forvar223} ?
          (reg228 != reg226) : (8'ha9)))));
      for (forvar237 = (1'h0); (forvar237 < (3'h4)); forvar237 = (forvar237 + (1'h1)))
        begin
          for (forvar238 = (1'h0); (forvar238 < (1'h1)); forvar238 = (forvar238 + (1'h1)))
            begin
              reg239 <= $unsigned((-$signed($unsigned((~^(8'ha4))))));
            end
          if ((-$unsigned(forvar238)))
            begin
              reg240 <= $unsigned((wire217 ?
                  ($signed(reg234) ?
                      {$unsigned(wire206),
                          (wire206 ?
                              reg236 : reg236)} : (|(forvar237 != wire208))) : {$signed({forvar223})}));
              reg241 = reg234;
              reg242 <= $unsigned("lZD14ok");
              reg243 <= forvar238[(3'h7):(3'h5)];
            end
          else
            begin
              reg240 <= wire217;
              reg241 <= reg213[(4'ha):(4'h9)];
            end
        end
      if ((($unsigned($signed(reg241)) ?
          (!(reg231[(2'h2):(1'h0)] ?
              reg226 : reg242[(1'h0):(1'h0)])) : reg219[(2'h2):(1'h0)]) ~^ (&($unsigned(forvar210) & ((!(8'had)) ?
          (forvar209 != reg240) : reg240[(3'h5):(1'h1)])))))
        begin
          if ({{(forvar238[(2'h3):(1'h1)] >= ((reg241 >= forvar237) << ((8'haf) || forvar223)))},
              forvar210[(5'h12):(4'hc)]})
            begin
              reg244 <= $unsigned((!((~(reg235 > reg215)) < (wire206 ?
                  (reg219 << reg234) : reg213[(3'h4):(2'h2)]))));
              reg245 = ($signed($unsigned(($unsigned(reg222) * wire208))) ?
                  $signed($signed({reg219})) : $signed({((!forvar210) >> forvar220[(3'h7):(3'h4)])}));
              reg246 <= $signed((reg226 ?
                  $signed($signed((reg239 ?
                      reg229 : forvar214))) : $signed($signed({forvar220,
                      reg245}))));
            end
          else
            begin
              reg244 = reg241[(4'ha):(1'h0)];
              reg245 = (reg234 ~^ (8'haa));
              reg246 <= $unsigned({((~^reg244) | {reg224}),
                  $unsigned(forvar223)});
            end
        end
      else
        begin
          if ("d")
            begin
              reg244 <= (~&$signed((+($signed(reg240) ?
                  forvar233[(3'h7):(3'h4)] : (reg236 >>> reg232)))));
              reg245 <= (^~(wire208 ^ $signed(wire208)));
              reg246 = reg227;
              reg247 = $unsigned((|((8'ha3) & reg224[(4'h8):(2'h2)])));
            end
          else
            begin
              reg244 = reg234[(1'h0):(1'h0)];
              reg245 = reg247;
              reg246 = {"yLmO1KmHJC55v3"};
              reg247 <= wire217;
              reg248 <= reg211;
            end
        end
      reg249 = (reg241 >> (reg232[(4'ha):(3'h6)] ?
          ($signed($signed(reg232)) ?
              reg242[(4'he):(4'h9)] : (7'h44)) : forvar209[(4'hc):(3'h6)]));
      reg250 = (!wire216[(1'h1):(1'h1)]);
    end
  assign wire251 = (-$unsigned(forvar210));
  assign wire252 = (8'hb4);
  assign wire253 = (|$unsigned({{forvar223[(4'h9):(3'h7)]}}));
  assign wire254 = ({wire217} ?
                       (({$unsigned(forvar223), $unsigned(reg243)} ?
                           ({reg242,
                               reg219} && $signed(reg248)) : reg234) == (8'hb6)) : (~^$unsigned(reg248)));
  always
    @(posedge clk) begin
      for (forvar255 = (1'h0); (forvar255 < (2'h3)); forvar255 = (forvar255 + (1'h1)))
        begin
          for (forvar256 = (1'h0); (forvar256 < (1'h1)); forvar256 = (forvar256 + (1'h1)))
            begin
              reg257 <= $signed(wire208[(3'h6):(2'h3)]);
              reg258 <= ($signed((reg244 && $unsigned((^~(8'hbb))))) >>> (($signed((~&reg218)) & $signed((~|forvar209))) ?
                  ((^~(8'hbf)) << ({wire253,
                      reg229} > (~^reg213))) : (+reg224)));
              reg259 <= {(reg235[(5'h10):(4'h9)] ? reg235 : $signed(reg227)),
                  forvar233[(2'h2):(2'h2)]};
              reg260 <= ($signed((~^$unsigned((forvar256 < reg225)))) ?
                  wire252 : reg230);
              reg261 = {({$unsigned($unsigned((7'h41))),
                      wire216} ~^ $signed({$unsigned(reg259)})),
                  (-(-(&$signed(forvar233))))};
            end
          if (reg225)
            begin
              reg262 <= $signed(forvar233);
              reg263 <= $unsigned(reg234);
              reg264 = (^reg219);
              reg265 = (8'hbc);
            end
          else
            begin
              reg262 <= (~^forvar210);
              reg263 <= reg249[(2'h2):(1'h0)];
              reg264 <= $unsigned(reg241);
              reg265 <= (-reg221[(2'h3):(2'h2)]);
            end
          for (forvar266 = (1'h0); (forvar266 < (1'h1)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 <= forvar220;
              reg268 = (~|wire252[(2'h3):(2'h3)]);
            end
          for (forvar269 = (1'h0); (forvar269 < (2'h3)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 <= $signed(reg264);
              reg271 <= (reg267 | reg259);
            end
        end
      for (forvar272 = (1'h0); (forvar272 < (1'h0)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 = $unsigned((reg260 && forvar237[(3'h4):(2'h3)]));
          reg274 <= (+(^(^$unsigned((-reg264)))));
          if (($unsigned(reg221) >>> reg273[(5'h12):(4'hb)]))
            begin
              reg275 <= $unsigned(reg257);
              reg276 = (reg244 < {(reg225[(2'h3):(1'h0)] ~^ ($signed(wire205) == (reg268 ?
                      reg222 : reg241))),
                  (reg222 == (8'hb6))});
            end
          else
            begin
              reg275 <= (reg265[(2'h2):(2'h2)] >>> $unsigned($signed($signed((reg212 ?
                  forvar266 : reg218)))));
            end
          for (forvar277 = (1'h0); (forvar277 < (2'h2)); forvar277 = (forvar277 + (1'h1)))
            begin
              reg278 <= forvar214;
            end
          for (forvar279 = (1'h0); (forvar279 < (1'h1)); forvar279 = (forvar279 + (1'h1)))
            begin
              reg280 = (~&(forvar214 ~^ $signed(reg260[(2'h3):(2'h3)])));
              reg281 <= (reg235 ?
                  ((("rSi" < (&(8'ha8))) ?
                          $signed(forvar266[(1'h0):(1'h0)]) : (reg211[(4'ha):(1'h0)] ?
                              $signed(wire252) : $signed(forvar256))) ?
                      $unsigned(($unsigned(reg218) > reg280)) : (~&((^reg228) ?
                          (reg259 != reg248) : reg261[(1'h1):(1'h1)]))) : reg267[(4'hb):(1'h0)]);
              reg282 <= ((reg215 ?
                      $signed(forvar237) : $signed(((reg225 == wire252) * $signed(reg221)))) ?
                  ({forvar233,
                      $signed($signed(wire251))} >> (((reg229 ~^ forvar266) || (reg234 + reg267)) ?
                      reg280[(1'h0):(1'h0)] : ($signed(reg270) ?
                          reg280[(1'h0):(1'h0)] : reg241))) : ($signed(reg270[(3'h4):(1'h0)]) ?
                      reg227 : $signed($unsigned((wire205 ?
                          wire206 : forvar237)))));
              reg283 = reg273[(4'hb):(4'hb)];
              reg284 = $signed(reg219[(4'hb):(3'h4)]);
            end
        end
    end
  assign wire285 = (!"");
  assign wire286 = $unsigned(((8'hbd) ?
                       (wire285[(2'h3):(2'h3)] || $signed(reg262[(4'he):(3'h6)])) : $signed((wire205[(1'h0):(1'h0)] == $unsigned(reg225)))));
  assign wire287 = $unsigned((({reg234, wire286[(5'h12):(4'hb)]} * reg239) ?
                       ((8'ha2) ?
                           (wire286 ?
                               (8'hab) : (reg257 != reg246)) : $unsigned((~|forvar272))) : $signed({$unsigned(reg250)})));
  assign wire288 = (((reg226[(2'h2):(1'h1)] <= $unsigned($unsigned(wire206))) != ($unsigned({forvar256}) ?
                           wire252 : ({reg228, reg270} ?
                               $signed(forvar220) : (~reg248)))) ?
                       (forvar266[(4'h8):(1'h1)] ?
                           (|reg248[(5'h10):(3'h5)]) : ($signed((reg271 ?
                                   reg219 : reg264)) ?
                               $signed(reg278) : (~|(reg257 ?
                                   (8'hbe) : reg267)))) : reg282);
  assign wire289 = (~|(reg275 + wire206));
  always
    @(posedge clk) begin
      if (reg240[(2'h3):(2'h2)])
        begin
          reg290 <= (reg232[(3'h5):(1'h0)] ?
              ($signed($unsigned((reg212 ?
                  reg231 : reg229))) >>> wire216) : (reg243 ?
                  ($unsigned((~|forvar279)) >= (^~reg265[(1'h1):(1'h0)])) : forvar255[(4'hc):(4'hb)]));
          for (forvar291 = (1'h0); (forvar291 < (2'h3)); forvar291 = (forvar291 + (1'h1)))
            begin
              reg292 = {$unsigned($unsigned(($unsigned(wire287) * reg274[(2'h2):(1'h0)])))};
              reg293 <= reg248[(5'h10):(4'h8)];
            end
          if ($signed($unsigned($unsigned(((forvar266 ?
              reg257 : wire288) >> ((8'hbb) ? forvar255 : reg264))))))
            begin
              reg294 <= {($signed((reg281 >>> forvar237)) <= {reg240[(2'h2):(1'h1)],
                      $unsigned($unsigned((8'hab)))}),
                  reg212[(1'h0):(1'h0)]};
              reg295 <= $unsigned(((($unsigned(reg226) ?
                      $signed(reg257) : wire251) ?
                  $signed((reg231 ^ reg225)) : $signed(wire285[(4'hc):(4'h8)])) <= $signed((8'ha3))));
              reg296 = (~($signed($unsigned((~|reg218))) || ((forvar220[(5'h10):(3'h6)] * {reg250,
                      wire217}) ?
                  (|((8'hbe) ^ wire207)) : reg236[(1'h1):(1'h1)])));
              reg297 <= ((&$signed(reg262[(4'he):(4'h9)])) >>> forvar223[(1'h1):(1'h0)]);
              reg298 <= {$unsigned((|(&(forvar238 <<< reg293)))),
                  {$unsigned($unsigned($unsigned(wire216))),
                      $unsigned($signed((reg265 >>> forvar238)))}};
            end
          else
            begin
              reg294 <= reg280[(2'h2):(1'h1)];
              reg295 <= wire205[(5'h12):(5'h10)];
              reg296 = (|(reg246[(3'h4):(2'h3)] ?
                  $unsigned(forvar269) : (^((reg267 ?
                      reg226 : reg290) != (reg219 >> reg241)))));
              reg297 <= wire288;
              reg298 <= $unsigned(reg245);
            end
          if ($unsigned(reg222[(4'h8):(4'h8)]))
            begin
              reg299 = {$unsigned(wire285), "wbMrMEY4FpLF8q3rT"};
              reg300 <= (~|$unsigned(wire288[(4'ha):(3'h6)]));
              reg301 <= reg282;
              reg302 <= $signed(reg259);
            end
          else
            begin
              reg299 = (8'hb8);
            end
        end
      else
        begin
          reg290 = $unsigned($signed({reg235[(3'h4):(2'h2)]}));
        end
    end
  always
    @(posedge clk) begin
      reg303 <= (wire289[(1'h0):(1'h0)] ?
          ((reg229 <<< (-(!reg226))) + $unsigned(reg301[(4'ha):(3'h5)])) : ($signed(reg218[(1'h0):(1'h0)]) <<< {"RhzxYnMXBw7Fo4T"}));
      reg304 = $signed($unsigned({(reg298 < reg293[(3'h7):(1'h0)]),
          reg247[(2'h2):(1'h0)]}));
      if ($signed({($signed(wire287) >> ($unsigned(reg234) ?
              $unsigned(reg229) : (^~wire205))),
          (((reg263 ? reg258 : (8'h9f)) ?
                  "e7aOh" : (reg244 ? reg219 : wire286)) ?
              $unsigned(((8'hb4) * reg225)) : "3iAapLsAYFg8KUmgbY")}))
        begin
          if (reg300[(1'h0):(1'h0)])
            begin
              reg305 = (($unsigned((forvar223 ?
                      (~&forvar214) : reg280[(2'h2):(1'h0)])) || ((^$signed((8'h9d))) ?
                      (^reg226) : (!{(8'hac)}))) ?
                  (7'h40) : $signed(reg301));
              reg306 <= (forvar223 && $unsigned($signed(reg258)));
              reg307 = ($unsigned((forvar269[(5'h14):(4'hc)] ?
                  {(reg232 ? (8'hac) : reg222),
                      (~reg232)} : ($unsigned(reg301) * $unsigned((8'had))))) ^ (((wire208[(3'h6):(1'h0)] ^ (reg224 >>> (7'h43))) >= ($unsigned(reg270) ?
                      wire206 : (reg271 ? reg262 : reg242))) ?
                  $unsigned($signed({reg267, forvar210})) : (8'ha1)));
              reg308 <= reg282;
              reg309 = reg265[(2'h2):(1'h0)];
            end
          else
            begin
              reg305 <= (reg257 ?
                  (({forvar291[(1'h1):(1'h0)]} ?
                      ((reg242 >= reg283) ^ reg290[(3'h6):(3'h4)]) : ($signed((8'hb7)) ?
                          $unsigned(reg304) : (reg248 & forvar269))) + $signed(((^reg295) ?
                      $signed(forvar256) : reg267))) : (reg212 ?
                      reg299 : reg260));
              reg306 = reg280;
              reg307 <= ((~^reg301[(3'h7):(3'h4)]) || forvar255[(3'h5):(2'h3)]);
              reg308 <= reg299[(4'hc):(2'h2)];
              reg309 <= $signed(reg248[(2'h3):(1'h1)]);
            end
        end
      else
        begin
          for (forvar305 = (1'h0); (forvar305 < (2'h3)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 = ($unsigned((+(8'h9f))) ?
                  (reg309[(3'h6):(3'h4)] == $unsigned(((~&reg239) ~^ reg240))) : ((reg259[(4'hb):(4'ha)] > "10weJbDklZ") <= reg212[(4'he):(4'hb)]));
              reg307 <= {$signed($unsigned($unsigned((reg234 | reg296)))),
                  $unsigned(reg218)};
              reg308 <= ((reg226 ?
                  $signed({$unsigned(reg239)}) : (!$unsigned(forvar237[(3'h7):(3'h7)]))) ~^ wire252);
            end
        end
      reg310 <= wire217;
      for (forvar311 = (1'h0); (forvar311 < (2'h3)); forvar311 = (forvar311 + (1'h1)))
        begin
          reg312 = $unsigned((reg244 >>> $unsigned(wire207[(4'h9):(3'h7)])));
          reg313 <= forvar279[(1'h1):(1'h1)];
          reg314 = (forvar209[(2'h2):(1'h0)] != $signed($unsigned(($signed(wire289) == $signed(reg308)))));
          reg315 <= ($unsigned({wire254,
                  ($signed(reg228) ? (+reg305) : $signed(reg247))}) ?
              (+$signed((8'hb2))) : ((^~{(wire254 ? forvar269 : reg297)}) ?
                  {(&reg294)} : (($unsigned(forvar237) || (wire286 + reg215)) > $signed((~reg261)))));
          for (forvar316 = (1'h0); (forvar316 < (1'h0)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 = (|"Z67FK");
              reg318 = wire254;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module27
#( parameter param168 = (((+(~&((8'ha3) ? (8'ha5) : (8'hb7)))) ? (~{((8'hb5) && (8'ha0)), ((8'h9e) <<< (8'hab))}) : ({((7'h42) >>> (7'h44))} | ({(8'ha0), (8'hae)} << (~^(8'hb8))))) ? ((^(((8'ha9) ? (8'hb7) : (7'h42)) ~^ (~^(8'ha6)))) ? ({((8'h9c) && (8'ha6))} ? ((~&(8'hbd)) && (~^(8'hbc))) : (((8'hb2) | (8'hb2)) ? (7'h40) : (&(8'haa)))) : {(((7'h44) * (8'ha6)) ? (~|(8'hb7)) : {(8'ha3)})}) : {(8'hbf)}) )
(y, clk, wire32, wire31, wire30, wire29, wire28);
  output wire [(32'h662):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire32;
  input wire [(4'h9):(1'h0)] wire31;
  input wire [(4'he):(1'h0)] wire30;
  input wire [(4'hd):(1'h0)] wire29;
  input wire signed [(3'h4):(1'h0)] wire28;
  wire signed [(3'h4):(1'h0)] wire167;
  wire [(3'h6):(1'h0)] wire166;
  reg [(5'h10):(1'h0)] reg165 = (1'h0);
  reg [(4'hb):(1'h0)] reg164 = (1'h0);
  reg [(5'h15):(1'h0)] reg163 = (1'h0);
  reg [(4'h9):(1'h0)] reg162 = (1'h0);
  reg [(2'h3):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg160 = (1'h0);
  reg [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar158 = (1'h0);
  reg [(3'h4):(1'h0)] reg157 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire156;
  wire [(4'h9):(1'h0)] wire155;
  wire signed [(5'h11):(1'h0)] wire154;
  reg signed [(5'h13):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg150 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg149 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar148 = (1'h0);
  reg [(3'h4):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] forvar144 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg145 = (1'h0);
  reg [(5'h13):(1'h0)] reg144 = (1'h0);
  reg [(5'h13):(1'h0)] reg135 = (1'h0);
  reg [(3'h4):(1'h0)] forvar133 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg143 = (1'h0);
  reg [(4'he):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg [(5'h13):(1'h0)] reg139 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg137 = (1'h0);
  reg [(4'ha):(1'h0)] reg136 = (1'h0);
  reg [(3'h5):(1'h0)] forvar135 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg134 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg133 = (1'h0);
  reg [(3'h7):(1'h0)] forvar132 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg129 = (1'h0);
  reg [(5'h13):(1'h0)] reg128 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar127 = (1'h0);
  reg [(3'h4):(1'h0)] reg126 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg125 = (1'h0);
  reg [(4'h9):(1'h0)] reg124 = (1'h0);
  reg [(4'hd):(1'h0)] reg123 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar121 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg119 = (1'h0);
  reg [(5'h13):(1'h0)] reg118 = (1'h0);
  reg [(4'hf):(1'h0)] forvar117 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg116 = (1'h0);
  reg [(2'h3):(1'h0)] reg115 = (1'h0);
  reg [(2'h2):(1'h0)] reg114 = (1'h0);
  reg [(4'hf):(1'h0)] forvar113 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg108 = (1'h0);
  reg [(2'h3):(1'h0)] reg107 = (1'h0);
  reg [(5'h11):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar105 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg104 = (1'h0);
  reg [(5'h15):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar101 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg100 = (1'h0);
  reg [(5'h11):(1'h0)] forvar99 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire98;
  reg signed [(4'h8):(1'h0)] reg97 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg96 = (1'h0);
  reg [(4'hc):(1'h0)] reg95 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg94 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg93 = (1'h0);
  reg [(5'h14):(1'h0)] forvar92 = (1'h0);
  reg [(2'h3):(1'h0)] reg91 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg90 = (1'h0);
  reg [(4'he):(1'h0)] reg89 = (1'h0);
  reg [(4'ha):(1'h0)] reg88 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg87 = (1'h0);
  reg [(5'h14):(1'h0)] forvar86 = (1'h0);
  reg [(3'h5):(1'h0)] reg85 = (1'h0);
  reg [(2'h2):(1'h0)] reg84 = (1'h0);
  reg [(4'hb):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg82 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg80 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar79 = (1'h0);
  reg [(4'he):(1'h0)] forvar78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg71 = (1'h0);
  reg [(5'h10):(1'h0)] forvar68 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar66 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg77 = (1'h0);
  reg [(4'h9):(1'h0)] reg76 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg75 = (1'h0);
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg [(4'h8):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg69 = (1'h0);
  reg [(2'h3):(1'h0)] reg68 = (1'h0);
  reg [(5'h13):(1'h0)] reg67 = (1'h0);
  reg [(5'h10):(1'h0)] reg66 = (1'h0);
  reg [(5'h12):(1'h0)] reg65 = (1'h0);
  reg [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg63 = (1'h0);
  reg [(4'he):(1'h0)] reg62 = (1'h0);
  reg [(4'ha):(1'h0)] reg61 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg60 = (1'h0);
  reg signed [(4'he):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar58 = (1'h0);
  reg [(5'h11):(1'h0)] reg57 = (1'h0);
  reg [(5'h11):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg55 = (1'h0);
  reg [(5'h13):(1'h0)] reg54 = (1'h0);
  reg [(4'ha):(1'h0)] reg53 = (1'h0);
  reg [(2'h3):(1'h0)] reg52 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg50 = (1'h0);
  reg [(4'hb):(1'h0)] reg49 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar48 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar45 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg44 = (1'h0);
  reg [(3'h4):(1'h0)] reg43 = (1'h0);
  reg signed [(4'he):(1'h0)] reg42 = (1'h0);
  reg signed [(4'he):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar40 = (1'h0);
  reg [(4'ha):(1'h0)] reg39 = (1'h0);
  reg [(5'h11):(1'h0)] forvar34 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg38 = (1'h0);
  reg [(4'h9):(1'h0)] reg37 = (1'h0);
  reg [(4'he):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg35 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg34 = (1'h0);
  wire [(3'h5):(1'h0)] wire33;
  assign y = {wire167,
                 wire166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 forvar158,
                 reg157,
                 wire156,
                 wire155,
                 wire154,
                 reg153,
                 reg152,
                 forvar151,
                 reg150,
                 reg149,
                 forvar148,
                 reg147,
                 reg146,
                 forvar144,
                 reg145,
                 reg144,
                 reg135,
                 forvar133,
                 reg132,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 reg133,
                 forvar132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 reg116,
                 reg115,
                 reg114,
                 forvar113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 forvar105,
                 reg104,
                 reg103,
                 reg102,
                 forvar101,
                 reg100,
                 forvar99,
                 wire98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 forvar92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 forvar86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 forvar79,
                 forvar78,
                 reg71,
                 forvar68,
                 forvar66,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 forvar71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 forvar58,
                 reg57,
                 reg48,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 forvar48,
                 reg47,
                 reg46,
                 forvar45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 forvar40,
                 reg39,
                 forvar34,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 wire33,
                 (1'h0)};
  assign wire33 = (wire28[(1'h0):(1'h0)] ?
                      (-wire31) : $signed($unsigned($unsigned(wire28))));
  always
    @(posedge clk) begin
      if ((($unsigned((+$unsigned(wire28))) && wire32[(3'h6):(3'h4)]) ?
          {(~(wire31 ?
                  $unsigned(wire31) : $signed(wire31)))} : wire28[(1'h1):(1'h0)]))
        begin
          if (wire28)
            begin
              reg34 <= (~|wire32);
              reg35 <= wire30;
              reg36 = $signed($signed(((&(~|wire30)) ?
                  (~&$signed(reg34)) : $signed({wire33, reg34}))));
              reg37 <= wire33[(3'h4):(2'h3)];
              reg38 <= (8'hb0);
            end
          else
            begin
              reg34 = ((reg38 ?
                      reg36[(3'h7):(3'h5)] : (~|{(reg37 ? wire28 : reg35),
                          {reg35}})) ?
                  {(^~$unsigned($unsigned(reg38)))} : $unsigned(reg36));
              reg35 <= $unsigned(reg36);
            end
        end
      else
        begin
          for (forvar34 = (1'h0); (forvar34 < (1'h0)); forvar34 = (forvar34 + (1'h1)))
            begin
              reg35 <= (reg37[(2'h2):(2'h2)] ?
                  $signed({($signed(reg34) ?
                          (^~(8'haf)) : (forvar34 > (8'hbb)))}) : reg37[(4'h9):(1'h0)]);
              reg36 = wire33[(3'h4):(1'h1)];
              reg37 = $signed((wire31[(1'h0):(1'h0)] ?
                  wire29 : (((wire29 ?
                      wire29 : reg34) & reg37) && ($unsigned(wire29) ?
                      (forvar34 && reg38) : reg34[(3'h5):(3'h4)]))));
              reg38 <= $signed($unsigned(wire29[(1'h0):(1'h0)]));
              reg39 = $unsigned(reg37[(1'h0):(1'h0)]);
            end
          for (forvar40 = (1'h0); (forvar40 < (1'h1)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 <= $unsigned($signed($unsigned("aVPCinoQRf0tPx")));
              reg42 <= ($unsigned(reg37[(2'h2):(1'h0)]) ?
                  (~(!(~(^reg36)))) : reg35[(3'h4):(2'h3)]);
              reg43 <= (8'h9d);
              reg44 <= (reg35 ?
                  (((~^reg41) ?
                          ("AQUCJcY" >> wire32[(3'h6):(2'h3)]) : (-(reg41 != wire28))) ?
                      $unsigned((reg34[(3'h5):(1'h0)] <= (~^(8'hbd)))) : (forvar34[(4'hf):(3'h5)] <= $unsigned(wire29))) : (reg36 - forvar40[(3'h7):(1'h1)]));
            end
        end
      if (wire32[(3'h5):(3'h4)])
        begin
          for (forvar45 = (1'h0); (forvar45 < (1'h1)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 = reg36[(4'hc):(4'h8)];
            end
          reg47 <= $signed(forvar34);
          for (forvar48 = (1'h0); (forvar48 < (2'h3)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 <= (~&(+$unsigned($unsigned((forvar48 & (8'ha2))))));
              reg50 <= $signed(reg46);
              reg51 = ((~forvar45) || reg36);
            end
          if ((8'hb1))
            begin
              reg52 <= (+($unsigned(reg37) ?
                  {$unsigned((reg42 ? reg38 : wire33))} : $signed(({(8'hb4),
                      wire28} ^~ (reg47 * wire28)))));
            end
          else
            begin
              reg52 <= $signed({$signed(reg44), $signed(reg51)});
              reg53 <= (($unsigned((~^(reg51 | (8'hb4)))) && "7lBoZS5ZNg9w3pkMm") ?
                  {"75D3YdbhNy"} : (8'hbe));
              reg54 = $signed((forvar34[(4'he):(4'hd)] ?
                  {(^wire29),
                      {(reg34 >> reg49),
                          reg51[(1'h0):(1'h0)]}} : $signed((wire30 ?
                      (wire29 ~^ reg43) : ((8'h9f) ? (8'ha3) : (8'ha0))))));
              reg55 = $signed(reg46[(3'h7):(2'h3)]);
              reg56 <= reg47[(2'h2):(1'h1)];
            end
        end
      else
        begin
          for (forvar45 = (1'h0); (forvar45 < (1'h0)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 <= (&reg41);
              reg47 <= $unsigned({reg56,
                  (reg55 ? reg39 : ((reg36 ? reg49 : (7'h42)) || forvar48))});
            end
          if (($unsigned("O2mGRG") + reg39))
            begin
              reg48 <= $signed({$signed("lrrTVUBul"),
                  ($signed($unsigned(reg51)) ?
                      ((reg36 ? reg54 : reg42) ?
                          (reg34 <<< reg39) : (^~wire33)) : reg36[(3'h6):(2'h3)])});
              reg49 <= {((~|(8'hb9)) & (|$signed((~|reg50))))};
              reg50 <= {($unsigned((reg47 && ((8'ha4) ?
                      reg47 : reg37))) | reg54)};
              reg51 = reg36;
            end
          else
            begin
              reg48 <= $signed($unsigned($unsigned({(reg46 ? reg53 : reg53)})));
            end
          reg52 <= reg50;
          if ($unsigned($signed(({$signed(reg49)} ?
              {$unsigned((8'h9f)), (8'h9f)} : forvar45))))
            begin
              reg53 <= wire28;
              reg54 <= ($unsigned(wire30) << ($signed(reg44) ?
                  (-$signed(reg49)) : $signed("kcA84VHsXzXPAhTmU2")));
            end
          else
            begin
              reg53 <= $unsigned(reg41);
              reg54 = forvar45;
              reg55 <= reg50;
              reg56 = $signed(forvar48[(3'h6):(1'h0)]);
              reg57 = ($unsigned((~^$unsigned((reg56 | reg39)))) == $unsigned($signed($unsigned($unsigned(reg42)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar58 = (1'h0); (forvar58 < (2'h2)); forvar58 = (forvar58 + (1'h1)))
        begin
          reg59 <= ($signed(wire29) ? reg54 : $unsigned((~(~^(|(8'hbe))))));
          reg60 = (((!(reg38 ? $signed(reg39) : "tsw8m")) >= (8'hb6)) ?
              forvar34 : $unsigned($unsigned($signed((~(8'ha8))))));
          if ($signed(($signed({(reg55 ? (7'h44) : reg35), (!reg53)}) ?
              ($unsigned({reg44}) ?
                  reg38 : $signed(reg34)) : $signed($signed("elJVdBhY3")))))
            begin
              reg61 = $signed((&((^(^(7'h42))) >> ((reg43 == wire30) ?
                  reg51 : $signed((8'ha1))))));
              reg62 = ($signed((forvar48[(3'h5):(3'h4)] ?
                      ((forvar34 ? reg60 : reg44) ?
                          $signed((7'h40)) : reg42[(4'hd):(4'hd)]) : $unsigned($unsigned(reg34)))) ?
                  $signed(reg35) : {((~&(!reg39)) ?
                          $unsigned(reg39) : (((8'haf) ?
                              reg42 : reg42) >>> reg54)),
                      reg43[(1'h0):(1'h0)]});
            end
          else
            begin
              reg61 <= ($signed($unsigned("MzM9awPu5l")) - forvar48);
              reg62 = $signed($unsigned((|$unsigned(reg49[(2'h3):(2'h3)]))));
              reg63 = (wire28 ?
                  ($signed(reg37[(3'h7):(3'h4)]) ?
                      $signed($signed($unsigned(reg46))) : $signed(forvar45)) : $signed(($unsigned($unsigned(reg57)) ?
                      (!(^wire33)) : wire28)));
            end
          reg64 <= reg37[(1'h1):(1'h1)];
        end
      if (reg54)
        begin
          reg65 <= $unsigned($unsigned((+$signed($signed(reg49)))));
          if ((|(~&$unsigned(reg43[(3'h4):(3'h4)]))))
            begin
              reg66 = reg52;
              reg67 <= forvar48;
              reg68 <= $unsigned(reg38);
              reg69 = ($unsigned(reg60) == wire33);
              reg70 <= {reg37[(1'h0):(1'h0)], $signed((8'h9d))};
            end
          else
            begin
              reg66 <= ((reg53[(3'h4):(2'h3)] >> wire32) ^ reg42[(2'h2):(2'h2)]);
              reg67 <= ($signed(((^(reg70 - reg38)) ?
                  (+((8'ha1) ^ reg41)) : $signed($signed(reg54)))) ~^ $signed(forvar40[(1'h0):(1'h0)]));
              reg68 = $unsigned(($unsigned(reg52[(1'h1):(1'h0)]) ?
                  $unsigned($signed((~^reg51))) : "Eskh7"));
            end
          for (forvar71 = (1'h0); (forvar71 < (2'h2)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 <= (reg57[(3'h5):(3'h5)] ?
                  reg61[(2'h2):(1'h0)] : {{reg41}});
              reg73 = $signed(reg38);
            end
          if ((reg63[(5'h11):(5'h11)] ?
              reg39[(3'h6):(1'h0)] : reg41[(2'h2):(1'h0)]))
            begin
              reg74 <= $unsigned(reg48[(4'h9):(3'h7)]);
              reg75 <= $signed(reg67[(5'h13):(4'hc)]);
              reg76 = (8'hab);
              reg77 = $unsigned(reg37);
            end
          else
            begin
              reg74 = (($unsigned({(!reg66),
                  (reg39 || reg62)}) ^ $unsigned(($signed(reg70) < $signed(reg62)))) << $unsigned($signed((~|(forvar58 | reg77)))));
            end
        end
      else
        begin
          reg65 = (($unsigned((forvar34[(4'he):(1'h0)] << "ePnnwPylUH08ek")) - reg38[(3'h7):(3'h4)]) > forvar34[(4'hf):(1'h1)]);
          for (forvar66 = (1'h0); (forvar66 < (3'h4)); forvar66 = (forvar66 + (1'h1)))
            begin
              reg67 <= ((^$signed(((reg56 - reg73) ?
                      (reg44 << reg74) : (forvar66 ? reg35 : reg59)))) ?
                  $unsigned((|({(8'ha8)} ?
                      "u81bGOLIRFROpAViO" : $unsigned(reg73)))) : $unsigned(reg34));
            end
          for (forvar68 = (1'h0); (forvar68 < (1'h0)); forvar68 = (forvar68 + (1'h1)))
            begin
              reg69 <= $unsigned($unsigned((reg59 ?
                  $signed(reg48[(2'h3):(2'h2)]) : wire28)));
              reg70 = forvar58;
              reg71 = ((reg73 ?
                      (reg67 ?
                          (-$signed(reg63)) : ($signed(reg67) - wire33)) : reg34[(2'h2):(1'h1)]) ?
                  reg66 : ({{(reg64 ? reg60 : (8'hbc))},
                      {wire29[(3'h5):(3'h5)],
                          $unsigned(wire28)}} < $signed((^(~|reg60)))));
              reg72 <= "0ffQgwurcT6BFvc";
              reg73 <= "IrpG2ScPThXtrZw4c";
            end
        end
      for (forvar78 = (1'h0); (forvar78 < (2'h3)); forvar78 = (forvar78 + (1'h1)))
        begin
          for (forvar79 = (1'h0); (forvar79 < (2'h2)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 <= (reg34[(2'h3):(2'h3)] ?
                  "iQz56TtMO3cTn1HDqmGa" : reg60[(2'h2):(1'h1)]);
              reg81 = (^{$unsigned({(reg55 - reg72), {reg34}}),
                  $unsigned($unsigned((reg59 ? (8'hbd) : (8'ha3))))});
              reg82 <= (|(reg48 ?
                  wire31[(1'h1):(1'h1)] : ((~|$unsigned(forvar40)) ?
                      $signed((forvar79 ? reg49 : reg48)) : ((reg44 ?
                              reg56 : reg55) ?
                          {(8'hbc)} : $unsigned(reg52)))));
              reg83 <= (reg52[(2'h2):(1'h1)] ?
                  $unsigned($signed(($signed((8'hbb)) ^ ((8'ha9) && reg56)))) : forvar40);
              reg84 = $signed($signed(((-(~^reg48)) ?
                  ((wire29 != (8'hac)) - $signed(reg66)) : {(reg83 && reg52),
                      $unsigned((8'haa))})));
            end
          reg85 = ({(forvar71 ? $unsigned((8'hae)) : $signed((8'hb5))),
              reg60[(2'h2):(1'h1)]} << (&$signed(reg70)));
          for (forvar86 = (1'h0); (forvar86 < (1'h1)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 <= {$signed(({(reg46 & reg81), (reg39 != reg37)} ?
                      ($unsigned(reg43) ^~ reg37[(3'h7):(1'h0)]) : (~|wire33)))};
              reg88 = reg35;
              reg89 <= $signed(((~&reg65[(2'h2):(2'h2)]) & wire29[(4'hb):(3'h5)]));
              reg90 <= wire30[(4'hb):(3'h6)];
            end
          if (reg36)
            begin
              reg91 = (reg46 | ((^($unsigned((8'hb8)) ?
                      ((8'hb2) ? reg64 : reg75) : reg66)) ?
                  (((8'hae) ? $unsigned((8'hb1)) : {reg66}) ?
                      reg55[(1'h1):(1'h0)] : ((reg71 ? reg61 : reg48) ?
                          reg53[(1'h0):(1'h0)] : (reg80 ?
                              wire28 : reg68))) : ((~^(~&reg37)) ?
                      (~(!reg77)) : forvar86)));
            end
          else
            begin
              reg91 <= ((($signed((reg39 | forvar68)) && ((reg83 + reg70) << (forvar45 ^ reg56))) != reg71[(2'h3):(2'h2)]) & $signed($signed((-"78O36HBKTx"))));
            end
          for (forvar92 = (1'h0); (forvar92 < (1'h0)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 <= forvar66;
              reg94 = reg54;
              reg95 = ($signed(reg85[(2'h3):(1'h1)]) ?
                  (("14ANXp930fq8d8mze" ?
                      (~&((8'ha0) + reg35)) : reg38[(4'he):(4'hd)]) ^ reg61[(1'h1):(1'h0)]) : reg52);
              reg96 = {(8'hac),
                  (^~(reg74 | ((reg95 >>> (8'hb4)) ?
                      $unsigned(reg49) : (reg81 << reg38))))};
              reg97 <= (($signed({$signed(reg73)}) ?
                      ((~^$unsigned(reg49)) || (7'h44)) : wire30) ?
                  $unsigned((reg38[(4'ha):(3'h7)] ^~ ({reg61, forvar86} ?
                      reg49 : reg83))) : $unsigned((^($signed(reg88) ?
                      $unsigned(reg91) : reg80[(1'h1):(1'h1)]))));
            end
        end
    end
  assign wire98 = (~^(+reg89[(3'h5):(1'h0)]));
  always
    @(posedge clk) begin
      for (forvar99 = (1'h0); (forvar99 < (2'h3)); forvar99 = (forvar99 + (1'h1)))
        begin
          reg100 = (($signed({(wire32 ?
                  reg35 : (8'hb9))}) && (~(7'h44))) ^~ ({reg68, (-(~^reg36))} ?
              forvar71[(2'h2):(2'h2)] : $unsigned((~^$signed(reg90)))));
          for (forvar101 = (1'h0); (forvar101 < (1'h1)); forvar101 = (forvar101 + (1'h1)))
            begin
              reg102 = reg53[(3'h6):(1'h1)];
              reg103 = ("RfdPymEUvyS" << {({{reg36, reg35}, (reg44 >>> reg75)} ?
                      $signed({forvar66, reg87}) : reg66),
                  ((+(wire32 < reg35)) ?
                      (~^(reg35 ?
                          (7'h44) : forvar79)) : (|reg66[(3'h5):(1'h0)]))});
              reg104 <= $signed($unsigned((!(^$signed(reg102)))));
            end
          for (forvar105 = (1'h0); (forvar105 < (2'h2)); forvar105 = (forvar105 + (1'h1)))
            begin
              reg106 <= ((~|$signed(((~^reg43) ?
                      (~reg59) : $unsigned(reg103)))) ?
                  $unsigned((reg70 ?
                      $unsigned(reg102[(4'ha):(2'h3)]) : $unsigned(reg74[(3'h6):(3'h5)]))) : reg67);
              reg107 <= $signed($unsigned($unsigned($unsigned(forvar66[(4'ha):(4'h9)]))));
              reg108 = reg71;
              reg109 <= {$unsigned(reg63[(5'h13):(4'hc)])};
              reg110 <= reg107[(2'h2):(2'h2)];
            end
          reg111 <= reg37[(1'h1):(1'h1)];
          reg112 = $unsigned((reg68 ?
              {"nSIxyq6qAMQURGVQ1xO"} : ($signed((reg102 ? reg88 : reg74)) ?
                  ((reg103 ^~ reg84) == $unsigned(wire33)) : forvar99[(3'h7):(2'h2)])));
        end
      for (forvar113 = (1'h0); (forvar113 < (2'h2)); forvar113 = (forvar113 + (1'h1)))
        begin
          if ({(reg109[(1'h0):(1'h0)] + ((+$unsigned(reg75)) ?
                  ($signed((8'ha8)) ? reg69 : reg42) : (~(reg109 ?
                      reg50 : reg37))))})
            begin
              reg114 = reg85;
              reg115 <= (|reg62[(1'h1):(1'h0)]);
              reg116 <= (8'hbd);
            end
          else
            begin
              reg114 <= {(~&($signed($unsigned(forvar113)) << (~&(~&forvar92)))),
                  wire29};
              reg115 <= reg41;
              reg116 <= $signed(reg51[(1'h1):(1'h1)]);
            end
          for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= (reg57[(3'h6):(3'h6)] ?
                  (^(-($unsigned(forvar113) - (8'hb4)))) : (reg35[(4'h9):(4'h8)] ?
                      (reg64 ?
                          ((-reg74) >>> {reg62,
                              reg55}) : $signed(((8'ha7) + forvar105))) : reg41));
              reg119 = $unsigned(reg88[(1'h1):(1'h0)]);
            end
          reg120 <= reg93;
          for (forvar121 = (1'h0); (forvar121 < (2'h3)); forvar121 = (forvar121 + (1'h1)))
            begin
              reg122 <= ((-wire33[(3'h5):(3'h5)]) ?
                  (($signed(((8'ha4) != forvar117)) ~^ $signed($unsigned(reg112))) ?
                      (^~(~|(reg34 || reg100))) : (|(&(~(8'h9c))))) : (-(+($unsigned(forvar117) ^ (-reg115)))));
              reg123 = (($signed(forvar68[(2'h3):(1'h1)]) < $unsigned((!forvar66))) >>> $unsigned(reg71[(4'ha):(2'h3)]));
              reg124 = (($unsigned({((8'ha0) ~^ reg66)}) || $unsigned($signed(wire29[(3'h6):(1'h0)]))) <= (~&(({reg123,
                      wire32} ?
                  (reg80 ?
                      (7'h44) : reg38) : (forvar86 >>> reg118)) ~^ (+(forvar86 ?
                  reg55 : (8'ha9))))));
              reg125 = ((wire32[(3'h4):(1'h1)] || ("u699Z96n" ?
                  $unsigned($unsigned(reg102)) : wire32)) - (^~(!(reg55 ?
                  {reg102, reg122} : (8'hb3)))));
              reg126 <= forvar121[(5'h11):(4'hf)];
            end
          for (forvar127 = (1'h0); (forvar127 < (2'h3)); forvar127 = (forvar127 + (1'h1)))
            begin
              reg128 <= reg110[(5'h10):(3'h7)];
              reg129 <= (-$unsigned(reg51[(1'h1):(1'h1)]));
              reg130 <= ($signed($signed((reg81 ~^ forvar117[(2'h3):(1'h0)]))) ?
                  (+$signed(($signed(forvar58) << $signed(reg83)))) : reg53[(2'h3):(1'h0)]);
              reg131 <= reg112;
            end
        end
    end
  always
    @(posedge clk) begin
      if ("7OrKqoB26usKouhPG7hR")
        begin
          for (forvar132 = (1'h0); (forvar132 < (3'h4)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= {((reg47[(1'h1):(1'h1)] ~^ $unsigned($signed(wire30))) ?
                      reg82 : (~reg115)),
                  $signed("81G4pc")};
            end
          reg134 = $signed(("YszhrM6vlSf3e" - (reg66 ?
              $unsigned(reg37) : $signed((8'hb6)))));
          for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= reg126[(3'h4):(1'h1)];
            end
          if ($unsigned(reg73))
            begin
              reg137 <= reg89[(4'he):(2'h2)];
              reg138 <= (~&(($unsigned(reg131) ?
                      $signed({reg35}) : wire28[(2'h3):(1'h1)]) ?
                  (((~|reg76) ? (&reg100) : ((8'hb2) != forvar117)) ?
                      $unsigned((forvar105 ? reg111 : reg120)) : ((+reg34) ?
                          (forvar40 ?
                              reg71 : (8'hb9)) : (forvar58 & reg110))) : reg88));
              reg139 <= $unsigned(((|$unsigned((reg55 && forvar105))) ?
                  (reg82[(5'h11):(3'h6)] ?
                      forvar101 : ((reg77 * reg34) < (~|reg46))) : $signed((8'hbc))));
              reg140 = reg136;
            end
          else
            begin
              reg137 <= reg139;
              reg138 <= $unsigned(($signed(reg118) ?
                  ($unsigned({reg93}) ?
                      $unsigned({reg80,
                          reg94}) : $signed(forvar117)) : reg106));
              reg139 <= $signed(reg41[(4'he):(4'he)]);
              reg140 = {reg72};
            end
          if ($unsigned(($unsigned(((^~reg139) ^~ $unsigned(reg140))) > $signed({reg139[(5'h13):(5'h13)]}))))
            begin
              reg141 <= $signed($signed((((reg76 ?
                  (8'hb7) : forvar117) > (8'ha7)) != reg74)));
              reg142 <= $signed(reg90);
            end
          else
            begin
              reg141 <= $signed(reg100);
              reg142 <= (~(!((~{reg72,
                  reg59}) || $unsigned($unsigned(reg67)))));
              reg143 <= reg41;
            end
        end
      else
        begin
          reg132 <= $unsigned(reg96[(2'h3):(1'h1)]);
          for (forvar133 = (1'h0); (forvar133 < (3'h4)); forvar133 = (forvar133 + (1'h1)))
            begin
              reg134 <= (($signed(({reg88} | $signed(wire30))) <= ((8'hb1) > forvar68[(4'he):(2'h2)])) ?
                  $signed($signed("vOkFfhJCRE32uI")) : $signed(reg108[(4'hd):(4'h8)]));
              reg135 <= "VYt2i1yHAI5E";
              reg136 <= $unsigned(((forvar121 ?
                      $signed((reg108 + reg94)) : reg84[(1'h1):(1'h0)]) ?
                  (7'h42) : "Yw2NnQ3hGunc50D"));
            end
          if (($unsigned(reg128) ?
              $unsigned($unsigned((reg122[(3'h5):(3'h5)] >>> $unsigned(reg66)))) : (((~|(forvar135 | reg109)) ?
                  ($signed(forvar92) > (|reg35)) : reg77) == ($signed($unsigned((7'h41))) == $signed((reg36 ?
                  reg39 : reg71))))))
            begin
              reg137 = (8'hb8);
            end
          else
            begin
              reg137 <= (8'ha9);
            end
          reg138 <= (~&reg131);
          reg139 = (reg83[(1'h0):(1'h0)] < $unsigned(forvar99[(4'hd):(4'hd)]));
        end
      if ({$unsigned($signed(reg49[(4'h9):(1'h0)]))})
        begin
          reg144 = {$signed($unsigned($signed((reg44 == reg47)))),
              (reg82[(2'h3):(2'h2)] ?
                  ($unsigned($unsigned(reg46)) & $signed(reg46[(2'h2):(2'h2)])) : {((~|forvar34) ?
                          reg106 : $signed(reg94))})};
          reg145 = (~{$signed(reg82[(1'h0):(1'h0)]),
              ($signed(reg51[(2'h2):(1'h0)]) == (^(reg50 ^~ reg46)))});
        end
      else
        begin
          for (forvar144 = (1'h0); (forvar144 < (2'h2)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 = reg75[(2'h3):(1'h1)];
              reg146 = $signed((reg114[(1'h1):(1'h1)] & "K2Bu"));
            end
          reg147 = $unsigned(($signed($unsigned(reg54)) ?
              $signed((forvar34 >= ((8'ha9) > forvar144))) : $unsigned("bSNhPM5")));
          for (forvar148 = (1'h0); (forvar148 < (2'h2)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 = reg111;
              reg150 = (("Vc1AKg5R4LJESA" != reg114) ?
                  ({"3s5bKepMp", "ytzYe"} ?
                      (({reg52,
                          (8'ha6)} <= reg42[(4'he):(3'h6)]) >>> forvar40[(3'h7):(3'h7)]) : (($unsigned(reg109) ?
                              $unsigned((8'hac)) : reg132[(2'h2):(2'h2)]) ?
                          $signed(forvar101) : {forvar144})) : (~&(forvar58 ^ (!((8'hbe) <= forvar45)))));
            end
          for (forvar151 = (1'h0); (forvar151 < (2'h2)); forvar151 = (forvar151 + (1'h1)))
            begin
              reg152 <= (($unsigned((reg97 ^~ $signed(reg67))) ^~ (~^((reg66 != reg46) != $signed(reg62)))) << $unsigned(reg68));
              reg153 = "8YpIrF9pCwTe3e4";
            end
        end
    end
  assign wire154 = ((8'h9c) ?
                       $unsigned(reg54) : $signed(($unsigned($unsigned(reg81)) ?
                           reg50 : $signed({reg77, reg46}))));
  assign wire155 = forvar71;
  assign wire156 = ($signed($signed({{reg35}})) ? reg50 : reg109);
  always
    @(posedge clk) begin
      reg157 <= $unsigned(($signed($unsigned((8'h9d))) != forvar92));
      for (forvar158 = (1'h0); (forvar158 < (1'h1)); forvar158 = (forvar158 + (1'h1)))
        begin
          reg159 <= $unsigned(($signed(reg71) << reg152[(4'h9):(3'h5)]));
          reg160 = $signed(reg122);
          if ((reg89[(4'hc):(1'h1)] ^~ {(~^reg124)}))
            begin
              reg161 = $unsigned($unsigned(($signed($signed((8'hba))) ?
                  (^~"1adtgqbK") : ($unsigned(forvar40) ?
                      ((7'h41) << reg44) : $signed(reg37)))));
              reg162 <= reg126[(1'h1):(1'h0)];
              reg163 <= reg109;
              reg164 <= ("K" || reg69);
              reg165 <= ($unsigned({({forvar78, reg95} && (8'hba))}) ?
                  (8'h9e) : $unsigned((reg143 - ($unsigned(wire29) <= $signed(wire33)))));
            end
          else
            begin
              reg161 <= "KMZANb4";
            end
        end
    end
  assign wire166 = (reg123 <= (forvar144[(3'h7):(2'h2)] ^ {"wk9Ck70kD1Q5E"}));
  assign wire167 = ($signed($signed(reg138)) || $unsigned($unsigned(((^~reg85) >= (~reg149)))));
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h106):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire4;
  input wire [(5'h10):(1'h0)] wire3;
  input wire signed [(4'h9):(1'h0)] wire2;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(5'h13):(1'h0)] wire0;
  wire signed [(5'h15):(1'h0)] wire164;
  wire [(4'h9):(1'h0)] wire162;
  wire signed [(5'h12):(1'h0)] wire28;
  wire signed [(4'hb):(1'h0)] wire18;
  wire [(4'hd):(1'h0)] wire17;
  wire signed [(5'h14):(1'h0)] wire16;
  wire signed [(2'h3):(1'h0)] wire15;
  wire [(5'h12):(1'h0)] wire14;
  wire [(5'h14):(1'h0)] wire13;
  wire [(4'h8):(1'h0)] wire12;
  wire signed [(4'hf):(1'h0)] wire11;
  wire signed [(5'h12):(1'h0)] wire10;
  wire signed [(5'h12):(1'h0)] wire9;
  wire [(5'h12):(1'h0)] wire8;
  wire signed [(4'h9):(1'h0)] wire7;
  wire signed [(5'h14):(1'h0)] wire160;
  reg signed [(4'hc):(1'h0)] reg6 = (1'h0);
  reg [(4'ha):(1'h0)] reg5 = (1'h0);
  assign y = {wire164,
                 wire162,
                 wire28,
                 wire18,
                 wire17,
                 wire16,
                 wire15,
                 wire14,
                 wire13,
                 wire12,
                 wire11,
                 wire10,
                 wire9,
                 wire8,
                 wire7,
                 wire160,
                 reg6,
                 reg5,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= $unsigned((wire4 ?
          wire0 : $signed((~(wire3 ? wire3 : (8'ha7))))));
      reg6 <= ((wire3[(4'hd):(3'h6)] * (8'hbd)) | $signed($signed(wire4[(5'h11):(3'h6)])));
    end
  assign wire7 = $unsigned((~&$signed(((reg6 ^~ reg6) ?
                     (wire3 ? (8'hb2) : wire2) : $unsigned(reg5)))));
  assign wire8 = wire1;
  assign wire9 = ($unsigned((wire0 + $unsigned({reg5}))) > $signed(($signed(wire0[(4'h9):(4'h8)]) ?
                     $signed((reg5 ~^ wire1)) : wire7)));
  assign wire10 = {$unsigned($unsigned((^wire3)))};
  assign wire11 = $unsigned((wire10[(4'hc):(4'h9)] ?
                      ({(~|reg6),
                          (~^wire1)} > $signed((wire9 & wire4))) : ($signed($unsigned(wire3)) ?
                          ((wire4 ? wire2 : wire9) ?
                              wire3 : reg5[(3'h7):(3'h4)]) : wire1[(4'hf):(2'h3)])));
  assign wire12 = wire11;
  assign wire13 = (+((~|reg6[(4'ha):(3'h7)]) ?
                      (wire8 ?
                          wire8 : $signed(((8'ha9) * wire10))) : ($signed(wire11) * $unsigned((wire4 ?
                          wire7 : wire1)))));
  assign wire14 = (wire12 ~^ $signed({(^(wire2 == wire9)), wire8}));
  assign wire15 = (~($signed(({wire4, wire12} ? (|wire8) : {wire7})) ?
                      $signed($unsigned(wire3[(4'hd):(1'h0)])) : (reg6 + wire8)));
  assign wire16 = ($signed(reg6[(1'h1):(1'h0)]) ?
                      (wire10 + $signed({(wire13 != wire12),
                          wire1[(1'h0):(1'h0)]})) : $signed((wire4[(4'hb):(2'h3)] ?
                          (^~wire3) : (+$signed(wire15)))));
  assign wire17 = $signed(((({wire4, wire15} + (reg5 ? wire4 : (8'h9c))) ?
                      (~^(wire9 ?
                          wire7 : wire10)) : ($unsigned(reg5) ^~ (wire7 && wire3))) > {((wire4 ?
                              wire8 : wire15) ?
                          wire2[(4'h8):(3'h4)] : ((8'h9e) ? wire16 : wire4)),
                      wire10}));
  assign wire18 = (wire14 ?
                      ((($unsigned(reg6) <<< (wire16 == wire16)) ?
                          $unsigned($unsigned((8'h9f))) : {((8'hb7) == (8'had)),
                              wire13}) || ((~&{wire1}) ?
                          reg5 : (8'hb8))) : $signed(wire8));
  module19 #() modinst29 (wire28, clk, reg5, wire1, wire18, wire0);
  module30 #() modinst161 (.wire31(wire28), .clk(clk), .y(wire160), .wire32(wire0), .wire33(wire14), .wire34(reg6));
  module30 #() modinst163 (wire162, clk, wire3, wire10, wire28, wire11);
  assign wire164 = ((wire9 <<< (((wire162 - wire14) <<< wire10) ?
                       (!(wire1 ?
                           wire1 : wire1)) : (&{reg6}))) | ({(wire2 >= wire9)} ?
                       wire11 : (+$unsigned(wire9[(4'h9):(3'h5)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module30  (y, clk, wire31, wire32, wire33, wire34);
  output wire [(32'h17a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire31;
  input wire signed [(5'h12):(1'h0)] wire32;
  input wire signed [(5'h12):(1'h0)] wire33;
  input wire signed [(4'ha):(1'h0)] wire34;
  wire [(4'hf):(1'h0)] wire159;
  wire [(3'h7):(1'h0)] wire158;
  wire signed [(5'h10):(1'h0)] wire157;
  wire signed [(5'h14):(1'h0)] wire35;
  wire signed [(2'h2):(1'h0)] wire64;
  wire [(5'h14):(1'h0)] wire66;
  wire [(3'h6):(1'h0)] wire71;
  wire [(5'h13):(1'h0)] wire91;
  wire signed [(3'h7):(1'h0)] wire93;
  wire signed [(3'h4):(1'h0)] wire94;
  wire [(4'hb):(1'h0)] wire95;
  wire [(4'hd):(1'h0)] wire96;
  wire [(3'h5):(1'h0)] wire97;
  wire signed [(5'h13):(1'h0)] wire98;
  wire [(4'h9):(1'h0)] wire108;
  wire signed [(4'he):(1'h0)] wire109;
  wire [(4'h9):(1'h0)] wire110;
  wire [(5'h13):(1'h0)] wire155;
  reg [(4'he):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg69 = (1'h0);
  reg [(3'h7):(1'h0)] reg68 = (1'h0);
  reg [(3'h6):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg102 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg105 = (1'h0);
  reg [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg107 = (1'h0);
  assign y = {wire159,
                 wire158,
                 wire157,
                 wire35,
                 wire64,
                 wire66,
                 wire71,
                 wire91,
                 wire93,
                 wire94,
                 wire95,
                 wire96,
                 wire97,
                 wire98,
                 wire108,
                 wire109,
                 wire110,
                 wire155,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 (1'h0)};
  assign wire35 = {wire32};
  module36 #() modinst65 (wire64, clk, wire32, wire35, wire34, wire33);
  assign wire66 = ((^$unsigned($signed((wire31 ? wire31 : wire33)))) ?
                      {($unsigned({wire32}) >> $signed((wire35 + (8'hb5))))} : wire31[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg67 <= $signed({wire64[(2'h2):(1'h1)]});
    end
  always
    @(posedge clk) begin
      reg68 <= $signed((|(8'hb2)));
      reg69 <= (({(8'hbe)} ?
              $unsigned((+$unsigned(wire66))) : $signed((~(wire64 != wire34)))) ?
          (wire64[(1'h1):(1'h0)] ?
              $signed($signed((^wire66))) : $unsigned(({wire64, (8'ha9)} ?
                  (wire33 << wire66) : (^~reg67)))) : ($unsigned(($unsigned((7'h43)) | (reg67 ?
                  wire34 : wire34))) ?
              ((^~(wire33 ?
                  reg68 : wire33)) + wire35) : wire35[(3'h4):(1'h1)]));
      reg70 <= (((($signed(reg68) ?
              {reg69, wire31} : $signed(wire33)) ^ (reg68 ?
              reg67 : (wire35 ?
                  (8'ha0) : wire32))) == (!(reg69[(2'h2):(2'h2)] & reg69))) ?
          ((8'ha7) ?
              ($unsigned(reg69[(3'h5):(2'h2)]) > ((wire66 ? wire34 : (8'hb2)) ?
                  $signed(wire32) : $unsigned(wire66))) : $signed($unsigned(wire34[(1'h1):(1'h0)]))) : {wire35[(1'h1):(1'h0)],
              wire31});
    end
  assign wire71 = (~$unsigned($unsigned(((^~(8'hb5)) ~^ (!reg68)))));
  module72 #() modinst92 (.wire75(reg69), .wire73(wire32), .y(wire91), .wire76(wire35), .wire77(wire66), .clk(clk), .wire74(wire31));
  assign wire93 = ({wire35} ?
                      {(($unsigned((8'hb9)) ?
                              wire31[(4'h9):(4'h9)] : (wire66 * (8'hbf))) || (~^wire35[(3'h7):(3'h4)]))} : $unsigned((({(8'hbf),
                          wire71} >>> wire91[(3'h5):(3'h5)]) + ((wire91 ?
                              reg67 : wire34) ?
                          wire66 : $signed(wire31)))));
  assign wire94 = reg67;
  assign wire95 = ((wire91 ~^ (($unsigned(wire94) ?
                              wire91[(4'hc):(2'h2)] : $signed(wire94)) ?
                          ($unsigned(wire34) ~^ $unsigned(wire34)) : ((reg67 ?
                                  wire71 : wire35) ?
                              wire71[(1'h1):(1'h0)] : {wire31}))) ?
                      (wire94 && $signed(wire32[(3'h4):(3'h4)])) : reg70);
  assign wire96 = wire31[(3'h6):(1'h1)];
  assign wire97 = {$signed((~wire96[(4'hc):(3'h6)])),
                      ({((8'hb7) ? $signed(wire71) : (^~wire31)), wire91} ?
                          $signed($unsigned(wire34[(1'h0):(1'h0)])) : ($unsigned(wire31) ?
                              $unsigned((8'hba)) : $signed((wire64 ?
                                  wire35 : wire64))))};
  assign wire98 = {{$signed(($unsigned(reg68) != $unsigned(wire31)))}};
  always
    @(posedge clk) begin
      if (((~|{reg70}) && (((!wire31[(2'h3):(1'h1)]) - wire35) ?
          $signed($signed(wire35)) : (!reg67[(2'h2):(1'h0)]))))
        begin
          reg99 <= ($signed($unsigned(reg68)) ?
              (((((8'ha0) && wire95) ?
                  wire35[(4'h8):(3'h7)] : reg69) & (wire96 > $signed(wire33))) == reg70[(4'ha):(3'h5)]) : $signed((|$signed((!wire94)))));
          reg100 <= wire64;
          reg101 <= reg100;
          reg102 <= wire33;
        end
      else
        begin
          if ((((reg67 > wire97[(1'h0):(1'h0)]) ?
                  $unsigned(((wire66 * wire93) || (|wire32))) : wire71) ?
              (wire31 ?
                  $signed((8'hb9)) : $signed($signed((wire33 ?
                      (7'h43) : reg99)))) : $signed(wire33[(4'h8):(3'h5)])))
            begin
              reg99 <= wire93;
              reg100 <= wire66;
              reg101 <= (wire71 ? $unsigned((8'h9c)) : wire98[(5'h13):(3'h6)]);
              reg102 <= $unsigned($signed((reg99[(2'h3):(1'h1)] & (^wire93[(3'h5):(3'h5)]))));
              reg103 <= {wire33,
                  $unsigned((wire33[(1'h1):(1'h1)] ?
                      ($unsigned((8'ha2)) || (!wire95)) : (wire95 ?
                          wire32[(3'h5):(3'h5)] : (wire93 <= reg69))))};
            end
          else
            begin
              reg99 <= $signed(({($unsigned(wire34) ?
                          (wire95 ? wire34 : wire71) : reg99)} ?
                  {$unsigned(reg68[(3'h7):(3'h4)])} : (!{{wire95, (8'ha8)}})));
              reg100 <= reg100;
            end
          if ($signed((((+{wire95}) * (^(wire96 == wire71))) + $unsigned(wire71[(3'h4):(3'h4)]))))
            begin
              reg104 <= $unsigned((8'ha1));
              reg105 <= wire97[(1'h0):(1'h0)];
            end
          else
            begin
              reg104 <= (wire33[(4'h9):(1'h0)] ? wire32 : reg102);
              reg105 <= reg69;
            end
        end
      if (wire96[(3'h6):(3'h4)])
        begin
          reg106 <= reg103;
        end
      else
        begin
          reg106 <= reg103[(1'h0):(1'h0)];
        end
      reg107 <= (reg69 ?
          (!(8'hab)) : $signed($unsigned(((^reg67) && wire97[(3'h4):(1'h0)]))));
    end
  assign wire108 = wire93[(3'h5):(1'h0)];
  assign wire109 = (wire71 << (&wire108));
  assign wire110 = {$unsigned($unsigned(((wire34 & wire98) ^~ (reg103 ?
                           wire98 : wire94))))};
  module111 #() modinst156 (.clk(clk), .wire112(reg106), .wire113(reg102), .wire115(wire33), .y(wire155), .wire114(reg69));
  assign wire157 = (~&(&$signed(reg99)));
  assign wire158 = reg99;
  assign wire159 = (+(8'hb2));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module19  (y, clk, wire23, wire22, wire21, wire20);
  output wire [(32'h23):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire23;
  input wire signed [(3'h5):(1'h0)] wire22;
  input wire [(3'h7):(1'h0)] wire21;
  input wire [(4'hd):(1'h0)] wire20;
  wire [(4'he):(1'h0)] wire27;
  wire signed [(2'h3):(1'h0)] wire26;
  wire signed [(4'he):(1'h0)] wire25;
  wire signed [(2'h3):(1'h0)] wire24;
  assign y = {wire27, wire26, wire25, wire24, (1'h0)};
  assign wire24 = $unsigned($unsigned((^~wire22)));
  assign wire25 = wire21[(2'h2):(1'h1)];
  assign wire26 = wire22[(2'h3):(1'h0)];
  assign wire27 = (({wire20[(4'hc):(4'ha)]} ?
                      ({(~|wire21),
                          {wire23,
                              wire21}} > ($signed(wire25) && (^~wire21))) : $unsigned(wire25[(4'h9):(1'h0)])) == ($signed({(&wire23)}) ?
                      ((|(8'haa)) ?
                          wire23[(4'ha):(2'h2)] : ((^~(8'hb4)) >= $unsigned(wire20))) : $signed($unsigned((wire20 ?
                          (8'hbc) : wire21)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module111
#(parameter param153 = ((~^(({(8'haa)} ? ((8'ha9) ? (8'ha3) : (7'h41)) : ((8'ha0) ? (8'hbb) : (8'ha1))) | (((7'h42) ~^ (8'hb9)) ? (!(8'haf)) : ((7'h41) >>> (8'hbf))))) ? (^~((^(~^(8'hba))) ? (((8'ha8) + (8'hab)) ? ((7'h44) * (8'hbb)) : (!(8'ha9))) : (((7'h40) > (8'hbe)) ? {(8'hbf)} : ((8'hbb) ^ (8'hb5))))) : ((^({(8'hbc)} ? ((8'h9f) ? (8'h9c) : (8'haf)) : ((8'haf) >= (8'hb3)))) ? (^~{(~&(8'h9d))}) : ((((8'ha1) ? (8'hbe) : (8'hb4)) ? (~|(8'hbc)) : ((8'ha8) || (8'haa))) ? ({(8'hb2), (8'hbd)} - {(8'hba), (8'hb1)}) : (~|(8'ha3))))), 
parameter param154 = {((((^(8'hae)) * (^~param153)) ? ((+(7'h44)) && (param153 ? param153 : param153)) : param153) ? {(param153 && (8'h9e))} : ((param153 ^ {param153}) ? (((8'haa) >= param153) + (~&param153)) : (param153 ? (8'hb9) : (+param153)))), (((+((8'haa) || (8'ha4))) <<< param153) - (~^{(param153 ~^ param153), (param153 ? param153 : param153)}))})
(y, clk, wire115, wire114, wire113, wire112);
  output wire [(32'h1ca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire115;
  input wire [(3'h7):(1'h0)] wire114;
  input wire signed [(5'h13):(1'h0)] wire113;
  input wire [(4'hb):(1'h0)] wire112;
  wire signed [(4'hd):(1'h0)] wire152;
  wire [(4'hd):(1'h0)] wire151;
  wire [(2'h3):(1'h0)] wire150;
  wire signed [(4'h8):(1'h0)] wire149;
  wire signed [(4'ha):(1'h0)] wire148;
  wire [(4'hd):(1'h0)] wire147;
  wire [(4'hf):(1'h0)] wire135;
  wire signed [(2'h3):(1'h0)] wire134;
  wire [(4'ha):(1'h0)] wire133;
  wire signed [(5'h14):(1'h0)] wire132;
  wire signed [(5'h15):(1'h0)] wire131;
  wire signed [(3'h7):(1'h0)] wire130;
  wire [(4'hc):(1'h0)] wire129;
  wire [(3'h4):(1'h0)] wire122;
  wire signed [(5'h14):(1'h0)] wire121;
  wire [(5'h13):(1'h0)] wire120;
  wire signed [(5'h11):(1'h0)] wire116;
  reg signed [(4'he):(1'h0)] reg146 = (1'h0);
  reg [(5'h14):(1'h0)] reg145 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg144 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg143 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg142 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg141 = (1'h0);
  reg [(3'h4):(1'h0)] reg140 = (1'h0);
  reg [(4'hc):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg127 = (1'h0);
  reg [(4'hb):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg123 = (1'h0);
  reg [(5'h12):(1'h0)] reg119 = (1'h0);
  reg [(4'h8):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg117 = (1'h0);
  assign y = {wire152,
                 wire151,
                 wire150,
                 wire149,
                 wire148,
                 wire147,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire131,
                 wire130,
                 wire129,
                 wire122,
                 wire121,
                 wire120,
                 wire116,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg119,
                 reg118,
                 reg117,
                 (1'h0)};
  assign wire116 = (8'haf);
  always
    @(posedge clk) begin
      reg117 <= $unsigned(wire112);
      reg118 <= wire114;
      reg119 <= $unsigned(((~^wire116[(1'h0):(1'h0)]) <<< $signed(((wire116 || wire116) ?
          $signed(wire114) : $unsigned(wire115)))));
    end
  assign wire120 = reg119;
  assign wire121 = wire112;
  assign wire122 = $signed((^~$unsigned(wire116[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      reg123 <= ($unsigned(wire120[(3'h5):(3'h5)]) ?
          reg119[(2'h2):(2'h2)] : ($signed(($unsigned(wire116) ?
                  $signed((8'h9d)) : (wire115 << wire115))) ?
              $signed($signed((reg117 >> (8'hae)))) : wire112[(3'h4):(2'h3)]));
      reg124 <= ((7'h40) >> $signed((wire116 ?
          ($unsigned(wire120) ?
              wire122 : wire120[(3'h4):(1'h0)]) : (^~(wire122 ?
              wire116 : wire115)))));
      reg125 <= ($unsigned($unsigned(((reg123 ?
          reg117 : wire121) ^~ wire122[(1'h1):(1'h1)]))) << (~^(8'hb7)));
      reg126 <= (+(+wire121));
      reg127 <= ($unsigned($unsigned({$signed(wire114),
          {(8'h9f), reg117}})) <<< $signed(($unsigned((wire113 ?
          (8'hbb) : (7'h43))) <= ($signed(reg118) - {reg117, (8'hae)}))));
    end
  always
    @(posedge clk) begin
      reg128 <= ((~|$signed(($unsigned(wire114) ^ $unsigned(reg127)))) ?
          $unsigned($signed(($signed((8'hbf)) ?
              (wire112 > wire120) : $signed(reg119)))) : ((^$signed($unsigned(reg119))) && reg117));
    end
  assign wire129 = $unsigned((~|{$signed(((8'hab) <= reg125))}));
  assign wire130 = {$signed(($signed(reg125) ? $unsigned((+reg127)) : reg125)),
                       wire122};
  assign wire131 = $signed($unsigned($signed(($unsigned(reg125) ?
                       (&(7'h43)) : reg127[(4'h9):(4'h9)]))));
  assign wire132 = (+$unsigned(((&{wire116}) + (+$unsigned(reg128)))));
  assign wire133 = wire120;
  assign wire134 = (~^{wire131});
  assign wire135 = $unsigned($signed((reg119[(3'h4):(2'h2)] ~^ reg123)));
  always
    @(posedge clk) begin
      reg136 <= (^$unsigned((|reg128[(4'hf):(3'h7)])));
      reg137 <= wire130[(3'h4):(2'h3)];
    end
  always
    @(posedge clk) begin
      if (wire134[(2'h3):(1'h0)])
        begin
          reg138 <= (({wire131[(4'hb):(3'h6)]} ?
              (((8'ha6) <<< $signed(wire129)) >> (~(wire134 ?
                  reg126 : reg137))) : reg137) << (+({$unsigned(reg119),
              (reg136 ? (8'hb0) : wire116)} <<< (8'ha6))));
          reg139 <= {$signed(reg127[(3'h7):(3'h7)])};
          reg140 <= (((^~{wire120, $signed(wire133)}) ?
              $unsigned($signed(wire133)) : $unsigned((-$signed(reg124)))) ~^ wire115[(5'h11):(3'h5)]);
        end
      else
        begin
          if ((8'hbc))
            begin
              reg138 <= {(wire130 ?
                      ({(~^wire131), (+reg138)} ?
                          $unsigned(wire130) : (reg140[(1'h1):(1'h1)] ?
                              (-wire121) : (~reg123))) : ((8'ha5) >>> $signed((+wire132))))};
              reg139 <= ((^~(reg136 < ((wire134 ? reg140 : reg124) ?
                  reg119 : (wire122 ?
                      wire132 : wire131)))) ~^ (!$signed($unsigned({reg124}))));
              reg140 <= {reg119};
              reg141 <= (^($signed($unsigned((reg118 ?
                  reg136 : wire130))) >> reg118));
            end
          else
            begin
              reg138 <= (reg137[(3'h6):(2'h3)] >= reg137);
              reg139 <= wire116;
            end
        end
      reg142 <= wire133[(4'ha):(3'h5)];
      if (wire113[(4'h8):(3'h7)])
        begin
          reg143 <= $unsigned($signed($unsigned({wire116})));
          reg144 <= wire133[(4'ha):(4'ha)];
          reg145 <= (reg128[(4'hb):(3'h7)] ?
              reg142[(3'h4):(1'h1)] : {{wire133}, reg128[(4'h8):(3'h5)]});
          reg146 <= $unsigned(reg125[(2'h2):(1'h0)]);
        end
      else
        begin
          reg143 <= wire120[(3'h7):(2'h3)];
          reg144 <= (^reg117);
          reg145 <= ({{$unsigned(wire115[(4'hf):(3'h5)])},
                  $signed(wire132[(3'h6):(2'h3)])} ?
              $unsigned($signed(($signed(wire120) > (wire115 != wire130)))) : (!$signed(wire116)));
          reg146 <= (wire116[(3'h4):(1'h1)] ?
              (~|(((wire115 ^~ wire135) - {(8'hb1)}) != $signed($signed((8'ha0))))) : (|(^~$signed({reg138,
                  wire129}))));
        end
    end
  assign wire147 = ((((~^$unsigned(reg126)) + (reg138[(4'h9):(4'h8)] ?
                           $unsigned(reg140) : (wire132 != reg136))) ?
                       (+(^~(reg144 ?
                           (8'h9c) : reg118))) : reg125[(3'h4):(1'h0)]) >> {wire122});
  assign wire148 = (~|(-$signed(reg126)));
  assign wire149 = $unsigned((($signed((reg136 == wire147)) ?
                           ((reg124 ?
                               wire112 : reg140) ^~ wire135[(4'hf):(4'he)]) : wire114) ?
                       reg136[(4'h8):(1'h1)] : ((+((8'h9e) ?
                               reg117 : wire133)) ?
                           (!$signed(reg125)) : reg137)));
  assign wire150 = reg139;
  assign wire151 = (wire131 ?
                       {(reg125[(1'h1):(1'h1)] ?
                               reg141 : (wire130[(2'h3):(2'h2)] >= $unsigned(wire120)))} : wire116[(3'h7):(3'h7)]);
  assign wire152 = reg119;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module72
#(parameter param89 = (((({(8'h9f)} ^~ (^(8'ha3))) - (((8'h9f) >= (8'haa)) ? (|(8'hb1)) : (!(8'hb3)))) ? (~|(^{(8'hac)})) : (+((~(8'hac)) + ((8'hb6) ? (8'ha2) : (8'ha4))))) - (({((8'hb5) << (8'hab)), ((8'ha3) && (8'haf))} ~^ (+((7'h42) ? (8'hab) : (8'h9e)))) ? (8'hb5) : {(~|((8'hb0) ? (8'ha1) : (8'hb4)))})), 
parameter param90 = param89)
(y, clk, wire77, wire76, wire75, wire74, wire73);
  output wire [(32'h6f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire77;
  input wire signed [(3'h5):(1'h0)] wire76;
  input wire [(4'h9):(1'h0)] wire75;
  input wire [(4'h9):(1'h0)] wire74;
  input wire [(3'h5):(1'h0)] wire73;
  wire [(4'hc):(1'h0)] wire88;
  wire [(5'h11):(1'h0)] wire87;
  wire [(4'hb):(1'h0)] wire86;
  wire [(4'h9):(1'h0)] wire85;
  wire signed [(2'h2):(1'h0)] wire84;
  wire [(4'hb):(1'h0)] wire83;
  wire [(4'hb):(1'h0)] wire82;
  wire signed [(2'h3):(1'h0)] wire78;
  reg signed [(4'h9):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg79 = (1'h0);
  assign y = {wire88,
                 wire87,
                 wire86,
                 wire85,
                 wire84,
                 wire83,
                 wire82,
                 wire78,
                 reg81,
                 reg80,
                 reg79,
                 (1'h0)};
  assign wire78 = wire76[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      reg79 <= wire78[(2'h3):(1'h1)];
      reg80 <= $unsigned((~&wire76));
      reg81 <= $signed($unsigned(wire74[(2'h2):(1'h1)]));
    end
  assign wire82 = $unsigned(reg79);
  assign wire83 = (+$signed(((^~(wire76 | wire82)) ?
                      wire74 : ((wire76 != reg81) < $signed(wire78)))));
  assign wire84 = ((-(~&$signed($unsigned(wire74)))) ? $signed(reg81) : wire77);
  assign wire85 = wire73;
  assign wire86 = wire84[(1'h1):(1'h0)];
  assign wire87 = {reg80, (~^wire78[(2'h3):(1'h0)])};
  assign wire88 = {wire86[(3'h5):(2'h2)],
                      ($signed(($signed((8'hbf)) ?
                              $unsigned(wire82) : $signed(wire82))) ?
                          wire73 : wire86[(2'h3):(2'h3)])};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module36
#(parameter param62 = ((8'hb2) >= (8'hb7)), 
parameter param63 = (8'hbc))
(y, clk, wire40, wire39, wire38, wire37);
  output wire [(32'hec):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire40;
  input wire [(5'h12):(1'h0)] wire39;
  input wire [(4'ha):(1'h0)] wire38;
  input wire signed [(4'ha):(1'h0)] wire37;
  wire [(4'hd):(1'h0)] wire59;
  wire signed [(4'h9):(1'h0)] wire53;
  wire signed [(4'h9):(1'h0)] wire52;
  wire signed [(5'h15):(1'h0)] wire51;
  wire [(4'hf):(1'h0)] wire50;
  wire [(4'hc):(1'h0)] wire49;
  wire [(3'h5):(1'h0)] wire48;
  wire signed [(5'h13):(1'h0)] wire47;
  wire [(3'h4):(1'h0)] wire46;
  wire signed [(4'hb):(1'h0)] wire45;
  wire [(4'hb):(1'h0)] wire44;
  wire signed [(4'ha):(1'h0)] wire43;
  wire [(3'h7):(1'h0)] wire42;
  wire [(3'h7):(1'h0)] wire41;
  reg [(5'h13):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg60 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg58 = (1'h0);
  reg [(5'h10):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(3'h7):(1'h0)] reg54 = (1'h0);
  assign y = {wire59,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 wire48,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 wire42,
                 wire41,
                 reg61,
                 reg60,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 (1'h0)};
  assign wire41 = {wire38};
  assign wire42 = wire40[(4'he):(4'h9)];
  assign wire43 = $unsigned(wire42);
  assign wire44 = (+(8'hbf));
  assign wire45 = (~&($unsigned(wire43[(4'h8):(4'h8)]) ?
                      (^~(wire40 ?
                          ((8'had) ? (8'hbe) : (8'h9d)) : (wire42 ?
                              (8'hb1) : wire42))) : {(8'ha9)}));
  assign wire46 = (^~$signed(wire41));
  assign wire47 = $signed({wire44[(4'hb):(4'hb)]});
  assign wire48 = (wire42[(1'h1):(1'h1)] | $unsigned(({$signed((8'h9f)),
                          (!wire44)} ?
                      $signed((wire38 ?
                          wire38 : (8'ha9))) : (wire46[(1'h1):(1'h0)] ?
                          wire40 : wire41[(3'h7):(3'h7)]))));
  assign wire49 = ($unsigned({$signed(wire46),
                      $unsigned((wire37 | wire48))}) >>> $signed(wire44));
  assign wire50 = ($unsigned($unsigned((wire49 ?
                      $signed(wire43) : wire38))) && ((~&(wire44 == {wire37,
                      wire37})) && wire43[(4'h8):(1'h0)]));
  assign wire51 = (~|wire48[(3'h4):(2'h3)]);
  assign wire52 = wire37;
  assign wire53 = wire50;
  always
    @(posedge clk) begin
      reg54 <= wire44;
      reg55 <= {$signed((^$signed((wire46 << wire51))))};
      reg56 <= (wire47[(3'h4):(3'h4)] ? wire46 : $unsigned(wire51));
      reg57 <= ($signed((!(^(^reg56)))) >> wire40[(4'he):(4'he)]);
      reg58 <= {wire41};
    end
  assign wire59 = ($signed(wire40[(3'h7):(1'h0)]) ?
                      (&(wire52 ?
                          (wire44 ?
                              $unsigned(wire43) : wire51) : wire45)) : wire42);
  always
    @(posedge clk) begin
      reg60 <= wire45;
      reg61 <= ((8'hb7) <= $signed((&wire41)));
    end
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param520 = (-(({(~^(7'h41)), ((8'h9e) ? (8'hb8) : (8'hb7))} ? ((~(8'hae)) - (~&(7'h43))) : (((8'had) == (8'hbe)) ? (!(8'h9f)) : (!(8'hb0)))) ? ((~^(~^(8'hb1))) ? (((8'ha8) << (8'hb9)) ? ((8'hbc) << (8'hb7)) : (~|(8'haa))) : (&(^(8'hb8)))) : ((((8'hb9) ? (7'h43) : (8'ha2)) && ((8'hb2) <= (7'h41))) ? {{(7'h42), (8'hb5)}} : ((~^(8'hb3)) < ((8'hb2) ? (8'ha4) : (8'ha7)))))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h3d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire0;
  input wire [(5'h11):(1'h0)] wire1;
  input wire signed [(4'ha):(1'h0)] wire2;
  input wire [(4'hb):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire4;
  wire signed [(5'h13):(1'h0)] wire5;
  wire signed [(2'h2):(1'h0)] wire6;
  wire signed [(5'h13):(1'h0)] wire7;
  wire signed [(5'h14):(1'h0)] wire518;
  assign y = {wire5, wire6, wire7, wire518, (1'h0)};
  assign wire5 = $signed($signed({("pvQQH" & $unsigned(wire4)), wire0}));
  assign wire6 = (wire0[(1'h0):(1'h0)] == $signed(wire5));
  assign wire7 = wire3;
  module8 #() modinst519 (wire518, clk, wire1, wire7, wire0, wire2, wire4);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module8
#(parameter param516 = ((((^((8'hbb) ? (8'h9f) : (8'h9e))) && (^~(^~(8'hbd)))) <= (!(((8'hbe) ? (8'hb7) : (8'h9c)) ? ((8'hac) ? (8'hb3) : (8'haa)) : (8'ha5)))) > ((~(((7'h42) ? (7'h40) : (8'hb7)) ? (8'hb7) : {(8'h9c)})) | ((((8'hbd) >>> (7'h44)) * (-(8'ha2))) || (^~((7'h41) >>> (8'ha5)))))), 
parameter param517 = (((8'h9e) < param516) && param516))
(y, clk, wire13, wire12, wire11, wire10, wire9);
  output wire [(32'h286):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire13;
  input wire [(5'h13):(1'h0)] wire12;
  input wire [(4'h9):(1'h0)] wire11;
  input wire [(4'ha):(1'h0)] wire10;
  input wire [(5'h11):(1'h0)] wire9;
  wire signed [(5'h13):(1'h0)] wire515;
  wire signed [(5'h15):(1'h0)] wire513;
  wire signed [(4'hc):(1'h0)] wire445;
  wire signed [(3'h6):(1'h0)] wire444;
  wire [(4'ha):(1'h0)] wire442;
  wire signed [(4'hc):(1'h0)] wire307;
  wire signed [(4'hc):(1'h0)] wire306;
  wire [(5'h13):(1'h0)] wire270;
  wire [(5'h11):(1'h0)] wire269;
  wire [(5'h13):(1'h0)] wire267;
  wire [(4'hb):(1'h0)] wire101;
  wire signed [(5'h15):(1'h0)] wire15;
  wire signed [(5'h13):(1'h0)] wire14;
  reg [(5'h11):(1'h0)] reg271 = (1'h0);
  reg [(4'h9):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg278 = (1'h0);
  reg [(4'hb):(1'h0)] reg279 = (1'h0);
  reg [(5'h14):(1'h0)] reg284 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg292 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg296 = (1'h0);
  reg [(5'h15):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg298 = (1'h0);
  reg [(4'ha):(1'h0)] reg300 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg302 = (1'h0);
  reg [(4'hc):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg305 = (1'h0);
  reg [(3'h4):(1'h0)] forvar303 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar301 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg299 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg295 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar294 = (1'h0);
  reg [(5'h10):(1'h0)] reg293 = (1'h0);
  reg [(2'h2):(1'h0)] reg291 = (1'h0);
  reg [(4'hd):(1'h0)] reg290 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar289 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar285 = (1'h0);
  reg [(5'h12):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg282 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar281 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar280 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg277 = (1'h0);
  reg [(2'h3):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar274 = (1'h0);
  reg [(4'hc):(1'h0)] forvar273 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg272 = (1'h0);
  reg [(2'h3):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg17 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg16 = (1'h0);
  assign y = {wire515,
                 wire513,
                 wire445,
                 wire444,
                 wire442,
                 wire307,
                 wire306,
                 wire270,
                 wire269,
                 wire267,
                 wire101,
                 wire15,
                 wire14,
                 reg271,
                 reg275,
                 reg278,
                 reg279,
                 reg284,
                 reg286,
                 reg287,
                 reg288,
                 reg292,
                 reg296,
                 reg297,
                 reg298,
                 reg300,
                 reg302,
                 reg304,
                 reg305,
                 forvar303,
                 forvar301,
                 reg299,
                 reg295,
                 forvar294,
                 reg293,
                 reg291,
                 reg290,
                 forvar289,
                 forvar285,
                 reg283,
                 reg282,
                 forvar281,
                 forvar280,
                 reg277,
                 reg276,
                 forvar274,
                 forvar273,
                 reg272,
                 reg18,
                 reg17,
                 reg16,
                 (1'h0)};
  assign wire14 = wire13;
  assign wire15 = $unsigned(wire11);
  always
    @(posedge clk) begin
      reg16 = $signed(((!$unsigned($unsigned(wire12))) << $unsigned({$unsigned(wire9)})));
      reg17 = $signed(wire13);
      reg18 = reg16[(3'h7):(3'h5)];
    end
  module19 #() modinst102 (.wire23(wire13), .wire21(wire12), .wire20(wire15), .wire22(wire9), .clk(clk), .y(wire101));
  module103 #() modinst268 (wire267, clk, wire15, wire13, wire14, wire101);
  assign wire269 = $signed($unsigned($unsigned(wire267)));
  assign wire270 = $signed(wire13[(3'h5):(2'h2)]);
  always
    @(posedge clk) begin
      reg271 <= ((&$unsigned(wire12[(3'h6):(3'h6)])) ?
          $unsigned((wire9 * $unsigned($signed(wire267)))) : (^~wire269));
      reg272 = $signed((~(wire10[(1'h0):(1'h0)] ?
          ({wire9} == (wire14 ?
              wire9 : wire270)) : $unsigned(wire9[(4'h9):(3'h6)]))));
      for (forvar273 = (1'h0); (forvar273 < (2'h2)); forvar273 = (forvar273 + (1'h1)))
        begin
          for (forvar274 = (1'h0); (forvar274 < (2'h2)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 <= wire15;
              reg276 = (8'ha0);
              reg277 = wire11[(4'h8):(2'h2)];
              reg278 <= (wire13[(2'h2):(1'h1)] * {{{((8'hb4) && (8'hb6))}}});
            end
        end
      reg279 <= wire11;
    end
  always
    @(posedge clk) begin
      for (forvar280 = (1'h0); (forvar280 < (1'h1)); forvar280 = (forvar280 + (1'h1)))
        begin
          for (forvar281 = (1'h0); (forvar281 < (1'h0)); forvar281 = (forvar281 + (1'h1)))
            begin
              reg282 = $signed($signed({($signed(wire9) ?
                      {wire9, wire14} : {forvar280})}));
              reg283 = ($signed((8'hb0)) ? wire101 : $unsigned(reg271));
              reg284 <= wire14[(4'he):(4'ha)];
            end
          for (forvar285 = (1'h0); (forvar285 < (1'h1)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 <= (reg271 ?
                  ((wire267 && $signed(wire11[(1'h0):(1'h0)])) ?
                      ("JtP3NlOxkppK" <= {(wire269 == reg282)}) : wire11[(4'h9):(3'h7)]) : reg275);
              reg287 <= $signed(wire12[(2'h2):(1'h1)]);
              reg288 <= wire12;
            end
          for (forvar289 = (1'h0); (forvar289 < (1'h1)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 = ({((^~{wire15}) | ((wire11 ? reg287 : wire14) ?
                          (wire9 > reg279) : (reg283 | wire10))),
                      {((wire267 <= wire14) ? (wire270 ^ wire270) : (8'hba))}} ?
                  {reg279,
                      $signed((8'hb1))} : ($unsigned(reg282) >> $unsigned(reg288)));
              reg291 = wire269;
              reg292 <= (wire269 + $unsigned($signed((^(wire10 <<< wire13)))));
              reg293 = wire13;
            end
          for (forvar294 = (1'h0); (forvar294 < (2'h3)); forvar294 = (forvar294 + (1'h1)))
            begin
              reg295 = wire9[(4'ha):(2'h3)];
            end
          if ($unsigned((wire12 ?
              forvar289 : (~|(wire10[(4'ha):(3'h6)] ?
                  (forvar280 ? (8'ha7) : reg283) : $unsigned(wire12))))))
            begin
              reg296 <= "v";
              reg297 <= (8'hbd);
              reg298 <= $signed((~|(7'h40)));
              reg299 = "ZB0a4OudHaTJwYgbayJr";
            end
          else
            begin
              reg296 <= $unsigned({wire9[(4'hf):(3'h7)]});
              reg297 <= ($signed((8'hbc)) ?
                  $unsigned((reg290[(1'h1):(1'h1)] ?
                      {((8'ha9) * reg291),
                          (forvar289 << reg283)} : reg295)) : reg296);
              reg298 <= $signed($signed(reg275[(3'h4):(2'h2)]));
              reg300 <= $signed(reg279);
            end
        end
      for (forvar301 = (1'h0); (forvar301 < (2'h2)); forvar301 = (forvar301 + (1'h1)))
        begin
          reg302 <= ((reg275[(2'h2):(1'h1)] ?
                  reg292[(2'h3):(2'h2)] : $signed((reg292 ^ $signed(reg286)))) ?
              reg282 : reg290[(3'h4):(1'h1)]);
          for (forvar303 = (1'h0); (forvar303 < (3'h4)); forvar303 = (forvar303 + (1'h1)))
            begin
              reg304 <= forvar285;
            end
        end
    end
  always
    @(posedge clk) begin
      reg305 <= $unsigned((8'hbb));
    end
  assign wire306 = $unsigned($unsigned((wire269[(2'h3):(1'h0)] <<< $unsigned(wire267[(3'h7):(2'h2)]))));
  assign wire307 = ($signed({reg292}) ?
                       wire9[(1'h0):(1'h0)] : (wire13[(3'h7):(1'h0)] || $signed(reg279)));
  module308 #() modinst443 (wire442, clk, wire270, reg297, wire10, reg287);
  assign wire444 = (~^{(-$signed((reg297 ? reg286 : reg278)))});
  assign wire445 = $unsigned((&(~|{(&wire270)})));
  module446 #() modinst514 (wire513, clk, reg271, wire269, wire267, reg300, reg279);
  assign wire515 = $unsigned("5B2VEygp70x");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module446
#(parameter param511 = {(({(~(8'hb5))} || (((8'hbd) && (8'hb7)) ? (!(8'h9f)) : ((8'ha6) ? (8'h9e) : (7'h42)))) << ((~|((8'had) ? (8'haf) : (8'ha7))) ? ({(8'h9e)} ? ((8'hbf) ? (8'hb1) : (8'hb6)) : {(8'hb4), (8'hb5)}) : (!((8'hb5) & (8'hb1))))), (+((((8'ha1) && (8'hbb)) ? {(8'ha3)} : (~^(7'h41))) ? ({(8'hbe), (8'hac)} >>> ((8'hb8) ^~ (8'hac))) : (^~((8'ha5) ? (8'hae) : (8'hbb)))))}, 
parameter param512 = (^~(((|param511) ? {(8'haf)} : (-((8'hb5) << param511))) && (((param511 >= param511) ^ {param511, param511}) ~^ ((param511 <<< param511) <= (^~(8'hae)))))))
(y, clk, wire451, wire450, wire449, wire448, wire447);
  output wire [(32'h302):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire451;
  input wire signed [(5'h11):(1'h0)] wire450;
  input wire signed [(3'h5):(1'h0)] wire449;
  input wire [(4'ha):(1'h0)] wire448;
  input wire [(4'hb):(1'h0)] wire447;
  wire [(2'h3):(1'h0)] wire470;
  wire [(4'hb):(1'h0)] wire469;
  wire [(5'h13):(1'h0)] wire468;
  wire [(5'h14):(1'h0)] wire467;
  wire signed [(4'hc):(1'h0)] wire466;
  wire [(3'h4):(1'h0)] wire465;
  wire [(3'h7):(1'h0)] wire464;
  wire [(4'ha):(1'h0)] wire463;
  wire signed [(5'h12):(1'h0)] wire462;
  reg signed [(4'hf):(1'h0)] reg510 = (1'h0);
  reg [(2'h2):(1'h0)] reg509 = (1'h0);
  reg [(3'h5):(1'h0)] reg508 = (1'h0);
  reg [(4'ha):(1'h0)] reg507 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg503 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg499 = (1'h0);
  reg [(4'hd):(1'h0)] reg498 = (1'h0);
  reg [(2'h2):(1'h0)] reg495 = (1'h0);
  reg [(2'h2):(1'h0)] reg491 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg489 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg487 = (1'h0);
  reg [(5'h15):(1'h0)] reg485 = (1'h0);
  reg [(5'h10):(1'h0)] reg484 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg481 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg479 = (1'h0);
  reg [(3'h6):(1'h0)] reg471 = (1'h0);
  reg [(4'he):(1'h0)] reg476 = (1'h0);
  reg [(3'h4):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg473 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg472 = (1'h0);
  reg [(3'h6):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg453 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg456 = (1'h0);
  reg [(3'h4):(1'h0)] reg455 = (1'h0);
  reg [(3'h5):(1'h0)] reg454 = (1'h0);
  reg [(4'hc):(1'h0)] reg452 = (1'h0);
  reg [(4'he):(1'h0)] reg506 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg505 = (1'h0);
  reg [(4'hd):(1'h0)] forvar504 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg502 = (1'h0);
  reg [(3'h6):(1'h0)] reg500 = (1'h0);
  reg [(5'h11):(1'h0)] reg497 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg496 = (1'h0);
  reg [(5'h13):(1'h0)] forvar493 = (1'h0);
  reg [(5'h11):(1'h0)] reg494 = (1'h0);
  reg [(5'h15):(1'h0)] reg493 = (1'h0);
  reg [(5'h13):(1'h0)] reg492 = (1'h0);
  reg [(5'h12):(1'h0)] reg488 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar486 = (1'h0);
  reg [(5'h14):(1'h0)] forvar481 = (1'h0);
  reg [(5'h13):(1'h0)] reg480 = (1'h0);
  reg [(4'h9):(1'h0)] reg483 = (1'h0);
  reg [(2'h2):(1'h0)] reg482 = (1'h0);
  reg [(5'h10):(1'h0)] forvar480 = (1'h0);
  reg [(5'h15):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar475 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg474 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar474 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar471 = (1'h0);
  reg [(4'ha):(1'h0)] reg460 = (1'h0);
  reg signed [(4'he):(1'h0)] reg459 = (1'h0);
  reg [(4'hf):(1'h0)] reg457 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar453 = (1'h0);
  assign y = {wire470,
                 wire469,
                 wire468,
                 wire467,
                 wire466,
                 wire465,
                 wire464,
                 wire463,
                 wire462,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg503,
                 reg501,
                 reg499,
                 reg498,
                 reg495,
                 reg491,
                 reg490,
                 reg489,
                 reg487,
                 reg485,
                 reg484,
                 reg481,
                 reg479,
                 reg471,
                 reg476,
                 reg475,
                 reg473,
                 reg472,
                 reg461,
                 reg458,
                 reg453,
                 reg456,
                 reg455,
                 reg454,
                 reg452,
                 reg506,
                 reg505,
                 forvar504,
                 reg502,
                 reg500,
                 reg497,
                 reg496,
                 forvar493,
                 reg494,
                 reg493,
                 reg492,
                 reg488,
                 forvar486,
                 forvar481,
                 reg480,
                 reg483,
                 reg482,
                 forvar480,
                 reg478,
                 reg477,
                 forvar475,
                 reg474,
                 forvar474,
                 forvar471,
                 reg460,
                 reg459,
                 reg457,
                 forvar453,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg452 <= (^~{((wire449[(3'h4):(2'h2)] ? (&wire450) : (^~wire449)) ?
              (wire451 ? {wire450, wire451} : {wire448}) : $signed(wire450))});
      if ((-{((wire447[(2'h3):(1'h0)] < {(8'h9d), wire448}) || wire450)}))
        begin
          for (forvar453 = (1'h0); (forvar453 < (1'h0)); forvar453 = (forvar453 + (1'h1)))
            begin
              reg454 <= $signed(wire448[(3'h7):(1'h1)]);
              reg455 <= $unsigned($unsigned($signed(($unsigned((8'hbe)) ^ (reg454 ?
                  (8'hb7) : reg452)))));
            end
          reg456 <= $unsigned($signed(wire447));
        end
      else
        begin
          if ($unsigned(wire448))
            begin
              reg453 <= $signed({wire448});
              reg457 = ($unsigned(wire448[(1'h0):(1'h0)]) | (($signed($signed(reg455)) ?
                  ((^(7'h43)) >> $signed(wire447)) : $signed(reg456[(2'h2):(1'h0)])) & (^~(wire450 ?
                  reg452[(2'h2):(1'h0)] : forvar453[(2'h2):(1'h1)]))));
              reg458 <= forvar453;
            end
          else
            begin
              reg457 = reg457[(4'h8):(1'h0)];
              reg458 <= {$unsigned({{forvar453[(1'h0):(1'h0)]},
                      ((wire451 ? reg457 : (8'haa)) ?
                          $unsigned(reg453) : {reg457})})};
              reg459 = $signed(wire451);
            end
          reg460 = reg453[(5'h10):(3'h5)];
        end
      reg461 <= ((8'hb8) - $signed(((&reg455) ?
          reg455[(3'h4):(2'h2)] : (!(reg454 ? reg453 : reg458)))));
    end
  assign wire462 = (-(($signed(reg456) || $signed(wire449)) | {((wire447 ?
                           wire451 : reg455) >= reg453)}));
  assign wire463 = (reg453 >>> ((!wire448[(2'h2):(1'h0)]) * reg461));
  assign wire464 = $signed($unsigned({(~&reg453), $unsigned((~reg456))}));
  assign wire465 = wire464;
  assign wire466 = ($signed((~|wire450)) ?
                       ($signed(($unsigned((8'haa)) ?
                               reg453[(5'h11):(2'h2)] : $unsigned((8'haf)))) ?
                           (~|(^~(^wire447))) : $unsigned($unsigned(((7'h42) ?
                               reg453 : reg452)))) : $unsigned($signed((8'ha8))));
  assign wire467 = $signed(reg455[(1'h1):(1'h1)]);
  assign wire468 = $unsigned((~^({(reg454 ~^ reg452)} ?
                       reg452[(4'h9):(4'h9)] : ($signed(wire464) ?
                           {reg461, reg456} : $signed(wire464)))));
  assign wire469 = (wire464 != wire465);
  assign wire470 = ($signed((reg461 < wire448)) & wire449);
  always
    @(posedge clk) begin
      if (((^{"nloOgd0UzA2M3rw0P77"}) ?
          $signed(($unsigned({wire449}) ?
              (reg455[(1'h1):(1'h1)] + "h") : (reg455 ^ wire451))) : ((((reg461 != reg454) ?
                  reg452[(3'h6):(3'h6)] : {reg461}) ?
              (wire448[(2'h3):(1'h1)] ~^ (wire469 ?
                  wire448 : reg456)) : (!$unsigned(wire470))) << wire462[(5'h12):(4'ha)])))
        begin
          for (forvar471 = (1'h0); (forvar471 < (2'h2)); forvar471 = (forvar471 + (1'h1)))
            begin
              reg472 <= (!$unsigned(($signed(wire467[(4'h9):(3'h4)]) == wire470[(2'h2):(1'h1)])));
              reg473 <= ($unsigned($signed((^forvar471[(3'h5):(2'h2)]))) * reg458[(5'h13):(5'h13)]);
            end
          for (forvar474 = (1'h0); (forvar474 < (1'h0)); forvar474 = (forvar474 + (1'h1)))
            begin
              reg475 <= $signed(reg472);
              reg476 <= forvar471;
            end
        end
      else
        begin
          if ($unsigned($signed(((~|(+(8'hb5))) ?
              $signed("yz5u8OJQy5v0ACh") : $signed({reg456})))))
            begin
              reg471 <= ((!(8'hbb)) ?
                  $signed((forvar471[(3'h5):(3'h5)] ?
                      (wire462[(3'h5):(1'h1)] ?
                          "k36dTNPP6E4ccIzhRt2" : wire462) : {(^reg473)})) : (reg453 ?
                      $unsigned(reg476[(4'hc):(2'h2)]) : wire467[(4'hc):(4'hb)]));
            end
          else
            begin
              reg471 <= (^~{$signed(($unsigned(reg454) || wire449[(3'h5):(1'h0)])),
                  reg454[(3'h4):(2'h3)]});
              reg474 = wire447[(3'h6):(3'h4)];
            end
          for (forvar475 = (1'h0); (forvar475 < (2'h3)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 <= (((~&($signed((8'h9c)) + (reg453 ?
                  reg452 : (8'ha3)))) + {$signed(wire449)}) >> (forvar475 ?
                  reg472[(4'hb):(1'h0)] : (wire449[(1'h1):(1'h0)] ?
                      $signed((wire469 > forvar475)) : $signed((~wire466)))));
              reg477 = (($unsigned($signed("CySUR8uXKn")) ?
                      $unsigned((!forvar475)) : (+(+reg474[(4'ha):(3'h6)]))) ?
                  forvar474 : ((~&wire462) ?
                      (wire465[(2'h2):(1'h0)] ?
                          ("HiVMVvY27pvF2Y" >> {reg453, reg472}) : ((^wire449) ?
                              reg461[(2'h3):(1'h0)] : reg453[(3'h6):(3'h6)])) : {(reg461[(1'h1):(1'h0)] ?
                              wire464[(2'h2):(1'h0)] : forvar471),
                          $signed((forvar471 || wire449))}));
              reg478 = ($signed((|$unsigned((^~reg475)))) ?
                  (8'haa) : ((~|$signed(((8'h9e) ? (8'hb4) : forvar475))) ?
                      $unsigned($signed("7h")) : {(^{reg477, forvar475}),
                          "47XVIU"}));
              reg479 <= (({{((8'hba) <= wire466),
                              (reg455 ? (8'ha5) : wire451)}} ?
                      forvar474 : wire449[(1'h1):(1'h0)]) ?
                  $signed(((~|{(8'hb9)}) ^ (-wire468))) : $signed($signed(($unsigned(wire467) >> (wire464 ?
                      reg474 : wire469)))));
            end
        end
      if (reg474)
        begin
          for (forvar480 = (1'h0); (forvar480 < (1'h1)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= (|((wire450[(1'h1):(1'h1)] > wire464[(3'h5):(1'h1)]) ?
                  (~$signed((wire465 ?
                      (8'hbd) : reg473))) : (~forvar475[(1'h1):(1'h0)])));
              reg482 = $unsigned((&wire467[(2'h3):(2'h2)]));
              reg483 = ($unsigned((((^~wire462) ?
                      (reg472 ? reg479 : reg479) : (&(8'h9d))) ?
                  $signed((wire449 ? reg456 : (8'hbc))) : ({forvar475} ?
                      $signed(wire450) : $signed(forvar480)))) | (($unsigned((wire469 <= reg455)) <= ((reg456 < wire450) <<< $unsigned(reg472))) ?
                  (!($unsigned(forvar474) ?
                      {reg461} : (reg452 > reg479))) : (8'ha1)));
            end
          reg484 <= ((+({(forvar475 - (8'ha8)),
                  (|reg471)} << (wire463 * (wire467 != reg472)))) ?
              ((~|wire449) ?
                  (+wire462) : $unsigned((wire467 & $unsigned((8'hb1))))) : wire451);
          reg485 <= (wire468 ?
              ($signed((^~$signed((8'hb3)))) ?
                  $unsigned($signed((reg481 ?
                      forvar471 : reg484))) : "RsEkbhcwrk7GCB") : (($signed({wire464,
                          reg477}) ?
                      reg472 : ((7'h40) + reg453)) ?
                  $signed(((~|forvar474) > reg453)) : $signed(($unsigned((8'hb3)) ?
                      $unsigned(wire463) : {wire467}))));
        end
      else
        begin
          reg480 = "IMIqO9OidL1u5";
          for (forvar481 = (1'h0); (forvar481 < (2'h3)); forvar481 = (forvar481 + (1'h1)))
            begin
              reg482 = "Lq6UD";
            end
        end
      for (forvar486 = (1'h0); (forvar486 < (2'h3)); forvar486 = (forvar486 + (1'h1)))
        begin
          if (((reg454[(1'h0):(1'h0)] ^ reg483[(4'h9):(3'h4)]) ?
              $signed($unsigned(($unsigned(reg452) >> reg455))) : $unsigned((((wire469 ?
                  reg461 : (8'hbb)) >= $signed((7'h44))) >>> (forvar474[(1'h0):(1'h0)] ?
                  ((8'h9d) * reg477) : $unsigned(forvar474))))))
            begin
              reg487 <= (8'ha4);
              reg488 = $unsigned(($signed($unsigned((~&forvar474))) ?
                  wire450[(4'ha):(3'h4)] : $signed(((+(8'hb9)) ?
                      (reg458 ? wire449 : wire464) : reg474[(4'h8):(1'h1)]))));
            end
          else
            begin
              reg487 <= ($unsigned(wire447[(2'h3):(2'h3)]) <= $unsigned(reg479));
            end
        end
      if ((~^reg485))
        begin
          reg489 <= ((((+reg487[(2'h3):(2'h2)]) & (((8'ha8) ?
                  reg488 : wire450) ?
              (reg456 ? reg480 : (8'haf)) : (reg485 ?
                  reg477 : wire468))) >>> {$unsigned(wire465[(3'h4):(2'h2)])}) | $unsigned(wire451[(3'h4):(2'h2)]));
          reg490 <= reg476[(4'h9):(1'h1)];
          if ((reg476[(4'h9):(1'h1)] > $unsigned(reg483)))
            begin
              reg491 <= $signed((reg481 ?
                  "W3RecloFKq5YVd" : $signed((reg479[(3'h4):(1'h1)] ?
                      reg474[(4'ha):(2'h2)] : $signed(wire466)))));
              reg492 = (reg454 ?
                  reg482 : ({reg473[(4'ha):(4'h9)]} ?
                      {$unsigned((reg454 > reg461))} : ($signed(wire447[(3'h7):(3'h7)]) ?
                          (reg482 ?
                              reg482[(2'h2):(1'h0)] : "xNW13yUtmHETMbisz") : reg456)));
              reg493 = (8'ha0);
              reg494 = "SXkN6";
            end
          else
            begin
              reg491 <= $signed($unsigned($unsigned((~^((8'ha0) ?
                  reg474 : reg491)))));
            end
        end
      else
        begin
          reg492 = (|$unsigned((forvar475[(1'h0):(1'h0)] && wire468)));
          for (forvar493 = (1'h0); (forvar493 < (3'h4)); forvar493 = (forvar493 + (1'h1)))
            begin
              reg494 = $signed($unsigned($unsigned((forvar493 == $unsigned(reg492)))));
              reg495 <= reg472;
              reg496 = $signed($unsigned((reg477[(3'h7):(3'h6)] & reg476[(4'hc):(2'h2)])));
              reg497 = ((~&(^~reg473[(1'h1):(1'h0)])) ?
                  reg452 : (!reg476[(3'h5):(2'h2)]));
              reg498 <= $signed(wire465);
            end
          if ($unsigned(wire467))
            begin
              reg499 <= $unsigned(wire468);
              reg500 = (reg461[(1'h1):(1'h0)] > $unsigned(reg479[(1'h1):(1'h0)]));
              reg501 <= {(8'hbc), "31HHrQz"};
              reg502 = (reg484[(4'ha):(1'h0)] ?
                  {forvar474,
                      (reg487[(3'h6):(2'h3)] == (~&reg485[(3'h5):(2'h3)]))} : reg456);
            end
          else
            begin
              reg499 <= (wire465[(1'h0):(1'h0)] >= forvar481);
              reg500 = $signed($signed(((8'h9c) ?
                  $signed((forvar474 ?
                      wire466 : reg489)) : wire470[(1'h1):(1'h0)])));
              reg501 <= (reg494[(1'h0):(1'h0)] - {(reg491 > forvar475[(1'h1):(1'h0)])});
              reg502 = $unsigned($unsigned($signed((reg497 == (reg461 >>> reg489)))));
              reg503 <= $unsigned(($signed($signed((~&reg487))) <<< (reg483 && ({reg484} ?
                  reg498[(3'h6):(1'h0)] : (!reg455)))));
            end
          for (forvar504 = (1'h0); (forvar504 < (2'h3)); forvar504 = (forvar504 + (1'h1)))
            begin
              reg505 = (reg499 ?
                  reg497[(3'h5):(2'h2)] : wire447[(3'h5):(1'h0)]);
              reg506 = ((|reg497[(4'hf):(4'hd)]) | $signed(wire448));
              reg507 <= ((8'hab) ? (8'hbe) : (^$unsigned((7'h42))));
              reg508 <= {((^forvar480[(3'h6):(1'h0)]) ?
                      ($signed(forvar493) ?
                          reg505[(3'h4):(1'h1)] : wire465[(1'h0):(1'h0)]) : (~|reg482)),
                  (($signed($unsigned(reg481)) * $unsigned($signed((8'hbb)))) ?
                      ($unsigned((wire463 ? reg487 : (8'ha8))) ?
                          (!(reg482 >> reg502)) : reg487) : (^{(wire462 == reg489),
                          $unsigned((8'hab))}))};
              reg509 <= reg497[(4'hb):(2'h3)];
            end
        end
      reg510 <= {reg475};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module308  (y, clk, wire312, wire311, wire310, wire309);
  output wire [(32'h61d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire312;
  input wire signed [(5'h15):(1'h0)] wire311;
  input wire signed [(3'h5):(1'h0)] wire310;
  input wire [(5'h15):(1'h0)] wire309;
  wire [(4'he):(1'h0)] wire415;
  wire [(3'h5):(1'h0)] wire389;
  wire signed [(4'he):(1'h0)] wire388;
  wire [(4'hd):(1'h0)] wire387;
  wire signed [(3'h4):(1'h0)] wire386;
  wire [(4'hf):(1'h0)] wire314;
  wire [(5'h13):(1'h0)] wire313;
  reg [(5'h15):(1'h0)] reg441 = (1'h0);
  reg signed [(4'he):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg436 = (1'h0);
  reg [(5'h10):(1'h0)] reg435 = (1'h0);
  reg [(2'h2):(1'h0)] reg433 = (1'h0);
  reg [(5'h12):(1'h0)] reg431 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg428 = (1'h0);
  reg [(4'h9):(1'h0)] reg420 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg414 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg413 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg411 = (1'h0);
  reg [(5'h13):(1'h0)] reg410 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg405 = (1'h0);
  reg [(4'he):(1'h0)] reg403 = (1'h0);
  reg [(5'h14):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg396 = (1'h0);
  reg [(4'hf):(1'h0)] reg395 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg394 = (1'h0);
  reg [(4'hf):(1'h0)] reg391 = (1'h0);
  reg [(4'h9):(1'h0)] reg385 = (1'h0);
  reg signed [(4'he):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg383 = (1'h0);
  reg [(2'h3):(1'h0)] reg380 = (1'h0);
  reg [(2'h3):(1'h0)] reg376 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg374 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg371 = (1'h0);
  reg [(5'h12):(1'h0)] reg369 = (1'h0);
  reg [(5'h12):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg365 = (1'h0);
  reg [(4'he):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg353 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg358 = (1'h0);
  reg [(5'h12):(1'h0)] reg357 = (1'h0);
  reg [(5'h13):(1'h0)] reg355 = (1'h0);
  reg [(2'h2):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg350 = (1'h0);
  reg [(4'h9):(1'h0)] reg348 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg347 = (1'h0);
  reg [(2'h3):(1'h0)] reg342 = (1'h0);
  reg [(5'h12):(1'h0)] reg339 = (1'h0);
  reg [(5'h12):(1'h0)] reg338 = (1'h0);
  reg [(4'h9):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg334 = (1'h0);
  reg [(3'h6):(1'h0)] reg332 = (1'h0);
  reg [(5'h13):(1'h0)] reg330 = (1'h0);
  reg [(5'h14):(1'h0)] reg328 = (1'h0);
  reg [(4'hd):(1'h0)] reg327 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg325 = (1'h0);
  reg [(3'h7):(1'h0)] reg324 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg323 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg319 = (1'h0);
  reg [(5'h12):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg439 = (1'h0);
  reg [(5'h12):(1'h0)] forvar438 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg434 = (1'h0);
  reg [(5'h15):(1'h0)] forvar432 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar430 = (1'h0);
  reg [(4'he):(1'h0)] reg429 = (1'h0);
  reg [(4'hb):(1'h0)] reg427 = (1'h0);
  reg [(4'h8):(1'h0)] reg426 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg425 = (1'h0);
  reg [(3'h7):(1'h0)] reg424 = (1'h0);
  reg [(5'h14):(1'h0)] forvar423 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar422 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg421 = (1'h0);
  reg [(4'hd):(1'h0)] reg419 = (1'h0);
  reg [(4'hb):(1'h0)] forvar418 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar417 = (1'h0);
  reg [(4'ha):(1'h0)] reg416 = (1'h0);
  reg [(4'h9):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg409 = (1'h0);
  reg [(4'h8):(1'h0)] reg408 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg407 = (1'h0);
  reg [(2'h2):(1'h0)] reg404 = (1'h0);
  reg [(3'h7):(1'h0)] reg402 = (1'h0);
  reg [(4'hf):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar397 = (1'h0);
  reg [(3'h6):(1'h0)] reg393 = (1'h0);
  reg signed [(4'he):(1'h0)] reg392 = (1'h0);
  reg [(5'h10):(1'h0)] forvar390 = (1'h0);
  reg [(3'h6):(1'h0)] reg382 = (1'h0);
  reg [(4'h9):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg379 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg377 = (1'h0);
  reg [(5'h14):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar367 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar366 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg349 = (1'h0);
  reg [(3'h4):(1'h0)] forvar348 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg361 = (1'h0);
  reg [(4'he):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar353 = (1'h0);
  reg [(4'ha):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar349 = (1'h0);
  reg [(5'h12):(1'h0)] forvar346 = (1'h0);
  reg signed [(4'he):(1'h0)] reg345 = (1'h0);
  reg [(3'h5):(1'h0)] reg344 = (1'h0);
  reg [(4'ha):(1'h0)] forvar343 = (1'h0);
  reg [(4'he):(1'h0)] forvar341 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg340 = (1'h0);
  reg [(4'he):(1'h0)] forvar336 = (1'h0);
  reg [(2'h2):(1'h0)] reg333 = (1'h0);
  reg [(5'h14):(1'h0)] forvar331 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg329 = (1'h0);
  reg [(2'h2):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg322 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar321 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg320 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg318 = (1'h0);
  reg [(5'h15):(1'h0)] reg317 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar316 = (1'h0);
  assign y = {wire415,
                 wire389,
                 wire388,
                 wire387,
                 wire386,
                 wire314,
                 wire313,
                 reg441,
                 reg440,
                 reg437,
                 reg436,
                 reg435,
                 reg433,
                 reg431,
                 reg428,
                 reg420,
                 reg414,
                 reg413,
                 reg411,
                 reg410,
                 reg406,
                 reg405,
                 reg403,
                 reg401,
                 reg400,
                 reg398,
                 reg396,
                 reg395,
                 reg394,
                 reg391,
                 reg385,
                 reg384,
                 reg383,
                 reg380,
                 reg376,
                 reg374,
                 reg373,
                 reg371,
                 reg369,
                 reg368,
                 reg365,
                 reg364,
                 reg353,
                 reg360,
                 reg358,
                 reg357,
                 reg355,
                 reg354,
                 reg352,
                 reg350,
                 reg348,
                 reg347,
                 reg342,
                 reg339,
                 reg338,
                 reg337,
                 reg335,
                 reg334,
                 reg332,
                 reg330,
                 reg328,
                 reg327,
                 reg325,
                 reg324,
                 reg323,
                 reg319,
                 reg315,
                 reg439,
                 forvar438,
                 reg434,
                 forvar432,
                 forvar430,
                 reg429,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 forvar423,
                 forvar422,
                 reg421,
                 reg419,
                 forvar418,
                 forvar417,
                 reg416,
                 reg412,
                 reg409,
                 reg408,
                 reg407,
                 reg404,
                 reg402,
                 reg399,
                 forvar397,
                 reg393,
                 reg392,
                 forvar390,
                 reg382,
                 reg381,
                 reg379,
                 forvar378,
                 reg377,
                 reg375,
                 reg372,
                 reg370,
                 forvar367,
                 forvar366,
                 reg363,
                 reg349,
                 forvar348,
                 reg362,
                 reg361,
                 reg359,
                 reg356,
                 forvar353,
                 reg351,
                 forvar349,
                 forvar346,
                 reg345,
                 reg344,
                 forvar343,
                 forvar341,
                 reg340,
                 forvar336,
                 reg333,
                 forvar331,
                 reg329,
                 reg326,
                 reg322,
                 forvar321,
                 reg320,
                 reg318,
                 reg317,
                 forvar316,
                 (1'h0)};
  assign wire313 = wire310;
  assign wire314 = $unsigned($unsigned(((~|$signed(wire310)) ?
                       ($unsigned(wire310) >= {wire310,
                           wire313}) : wire313[(4'h9):(1'h0)])));
  always
    @(posedge clk) begin
      reg315 <= (-(8'haa));
      for (forvar316 = (1'h0); (forvar316 < (1'h1)); forvar316 = (forvar316 + (1'h1)))
        begin
          if (((^forvar316[(1'h1):(1'h0)]) >= $signed(((&wire314[(4'hd):(3'h4)]) >>> $signed($signed(reg315))))))
            begin
              reg317 = wire311[(5'h15):(4'hf)];
              reg318 = ((&wire310[(1'h0):(1'h0)]) ~^ reg315[(1'h1):(1'h1)]);
              reg319 <= $signed(($signed($unsigned($unsigned(forvar316))) ^~ reg317[(4'he):(4'hb)]));
              reg320 = (^reg318);
            end
          else
            begin
              reg319 <= wire311[(4'he):(1'h0)];
              reg320 = {(forvar316[(2'h2):(1'h0)] ?
                      (reg317[(1'h0):(1'h0)] && $signed((wire311 << wire309))) : wire309),
                  (wire311[(4'h9):(3'h6)] ?
                      $unsigned(reg318[(3'h5):(3'h5)]) : wire309)};
            end
          for (forvar321 = (1'h0); (forvar321 < (1'h0)); forvar321 = (forvar321 + (1'h1)))
            begin
              reg322 = (+($signed(reg320[(1'h1):(1'h0)]) ?
                  $unsigned(($signed(reg320) ?
                      ((8'hba) ?
                          wire311 : forvar321) : (wire311 <= wire313))) : reg320));
              reg323 <= ($unsigned((reg322[(2'h2):(1'h0)] & wire314[(1'h0):(1'h0)])) > wire312);
              reg324 <= (wire312[(3'h7):(3'h4)] ?
                  (reg322 ?
                      wire312[(3'h4):(1'h0)] : $signed({{(7'h42)}})) : forvar316);
              reg325 <= reg318;
              reg326 = ({(($signed(forvar316) * $unsigned(forvar316)) ?
                      ((reg317 ? (8'hb1) : reg319) ?
                          (reg323 != wire312) : reg315[(4'h9):(3'h6)]) : wire311),
                  (8'haf)} | $signed($unsigned((^""))));
            end
        end
      if (forvar321)
        begin
          reg327 <= (-(($signed((~&reg323)) << $unsigned($signed((8'ha4)))) & ((reg323 != $unsigned(reg317)) ?
              ({reg315} ? $unsigned(reg322) : reg322) : wire311)));
          if ("TMBVLt6UoQcEw2D4TalT")
            begin
              reg328 <= $unsigned((reg325 >>> (8'hab)));
              reg329 = (^((-$unsigned({wire311,
                  (8'hb6)})) ~^ {((^~reg320) ~^ (~&reg317)),
                  {wire314[(3'h5):(2'h2)]}}));
            end
          else
            begin
              reg328 <= (((!$signed((reg326 <= reg323))) * $signed(reg328)) != forvar316[(1'h0):(1'h0)]);
              reg329 = ("q7vdikzf29Aw" ~^ {reg329[(5'h10):(4'h9)],
                  reg315[(4'hd):(1'h1)]});
            end
          reg330 <= (~|$unsigned({(^~$signed(reg326))}));
          for (forvar331 = (1'h0); (forvar331 < (3'h4)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 <= (wire309[(4'hf):(3'h4)] ?
                  ((^~wire310) ?
                      reg324 : (+$signed(forvar321))) : $signed((-((^~forvar331) << (reg320 ?
                      (8'hb0) : reg320)))));
              reg333 = wire313[(5'h11):(3'h6)];
              reg334 <= ($signed(reg329) ?
                  reg324 : (reg320[(2'h3):(1'h1)] == $unsigned((&reg319[(4'ha):(4'ha)]))));
              reg335 <= {$signed(wire314)};
            end
        end
      else
        begin
          reg327 <= (7'h42);
        end
      for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
        begin
          reg337 <= reg320[(3'h4):(1'h0)];
          reg338 <= reg330[(4'he):(4'h8)];
          reg339 <= (reg319[(3'h7):(3'h7)] && (reg330[(4'hb):(3'h7)] + $unsigned($unsigned(wire313))));
          reg340 = ($signed((~&(^$signed(reg328)))) || $unsigned($unsigned({(8'ha8)})));
        end
    end
  always
    @(posedge clk) begin
      for (forvar341 = (1'h0); (forvar341 < (1'h1)); forvar341 = (forvar341 + (1'h1)))
        begin
          reg342 <= (~&(((^~((8'h9e) <<< (8'ha2))) | reg327) | (reg338[(4'h8):(2'h3)] ?
              {reg324, $signed(wire314)} : $signed("1qOVkIdEJHbP1AUA"))));
          for (forvar343 = (1'h0); (forvar343 < (1'h0)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 = reg338[(1'h0):(1'h0)];
              reg345 = reg339;
            end
          for (forvar346 = (1'h0); (forvar346 < (2'h3)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 <= $unsigned("IvDY1n1T");
            end
        end
      if ($signed(((!$signed(reg315[(4'he):(1'h1)])) ?
          (^~{forvar341[(3'h4):(1'h1)]}) : ((8'ha0) ?
              $unsigned((8'hb3)) : (reg334 << $unsigned(wire314))))))
        begin
          reg348 <= reg339[(4'he):(3'h6)];
          for (forvar349 = (1'h0); (forvar349 < (2'h2)); forvar349 = (forvar349 + (1'h1)))
            begin
              reg350 <= $signed((~&$unsigned((~(reg324 | (8'hba))))));
              reg351 = {(~$signed(reg342[(1'h0):(1'h0)]))};
            end
          reg352 <= $unsigned((~|(((8'h9d) ?
              (~|reg350) : $unsigned(wire310)) * $signed($signed(reg351)))));
          for (forvar353 = (1'h0); (forvar353 < (1'h1)); forvar353 = (forvar353 + (1'h1)))
            begin
              reg354 <= $signed(reg324[(2'h2):(1'h0)]);
              reg355 <= reg348;
              reg356 = ($unsigned(("tNai6KVr4" ?
                  "" : reg337)) * $signed($unsigned($unsigned({(8'ha4),
                  reg350}))));
            end
          if (($unsigned(reg352) ?
              (^~reg325[(2'h3):(2'h3)]) : ((reg348 ?
                  ((8'haa) - "hPPVgqRKKyYBvJ5fu") : $unsigned((|reg351))) == reg350[(3'h6):(2'h3)])))
            begin
              reg357 <= reg324;
              reg358 <= (+(reg351 ?
                  $signed((^(forvar353 ^~ reg354))) : (wire314 ?
                      ((reg357 == wire314) ?
                          reg356 : reg344[(3'h4):(3'h4)]) : $unsigned($unsigned(reg325)))));
            end
          else
            begin
              reg359 = ((reg324[(3'h7):(1'h1)] ^ $unsigned($unsigned((7'h43)))) ?
                  reg327[(4'hc):(3'h6)] : (($signed((~^forvar346)) ?
                      reg327 : ((-reg345) >> {reg323,
                          reg332})) >= "2wwtSG7UDub8h1MoU0"));
              reg360 <= $signed((({"V6y"} | $signed((~^(8'hbd)))) ?
                  $signed({((8'h9e) ?
                          wire312 : (8'hb4))}) : reg328[(5'h13):(4'hc)]));
              reg361 = wire314;
              reg362 = {reg348, $signed($signed(reg345))};
            end
        end
      else
        begin
          for (forvar348 = (1'h0); (forvar348 < (1'h0)); forvar348 = (forvar348 + (1'h1)))
            begin
              reg349 = reg358[(3'h4):(2'h2)];
              reg351 = (~&(reg358[(5'h10):(4'hc)] ?
                  reg339 : wire311[(4'hc):(4'hc)]));
              reg352 <= $unsigned($signed($signed((reg328 <= reg328[(4'hd):(2'h3)]))));
              reg353 <= (($signed(((~&reg349) ?
                  (+reg348) : $unsigned(reg355))) ^~ $signed((8'ha4))) ~^ $unsigned((~|$signed(((8'ha0) ^ reg347)))));
              reg356 = (~|"UopDUUVgdbGizkDezu");
            end
          reg359 = $signed((~&(($unsigned(reg361) <= (^reg356)) <<< reg361)));
          reg360 <= $signed(($signed((~&reg355[(3'h6):(3'h6)])) ^~ $signed(reg362[(4'h8):(2'h2)])));
          if (reg355[(1'h1):(1'h0)])
            begin
              reg361 = reg354;
              reg362 = (8'hbe);
            end
          else
            begin
              reg361 = $unsigned($unsigned({$unsigned(((8'ha1) != reg351))}));
            end
          reg363 = $signed((|(|((^(8'had)) + wire312[(1'h1):(1'h1)]))));
        end
      reg364 <= ((reg361 ?
              ($unsigned((!reg330)) - ((8'ha7) >>> (-wire309))) : ($signed($unsigned(forvar346)) | $unsigned("tsPCL"))) ?
          ((^{$unsigned(reg358)}) + reg338) : $unsigned((-((reg332 ?
                  wire310 : (8'ha7)) ?
              (+(8'h9d)) : {reg356}))));
      reg365 <= (reg344 ?
          $signed(wire312[(2'h3):(2'h2)]) : reg356[(5'h11):(3'h7)]);
      for (forvar366 = (1'h0); (forvar366 < (1'h1)); forvar366 = (forvar366 + (1'h1)))
        begin
          for (forvar367 = (1'h0); (forvar367 < (1'h1)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 <= (8'hb0);
              reg369 <= $unsigned(reg347);
              reg370 = $signed($unsigned((~&$unsigned($signed(reg328)))));
            end
          if ($signed(reg355))
            begin
              reg371 <= (7'h41);
              reg372 = (+(^~reg358[(4'hb):(4'ha)]));
            end
          else
            begin
              reg371 <= ($unsigned($signed(($unsigned(reg360) ?
                  wire314 : reg359))) >= $unsigned($signed(reg351[(3'h4):(2'h3)])));
              reg373 <= (!{(+reg364)});
              reg374 <= ($signed(reg353[(4'h8):(3'h7)]) - (^~(($signed(reg359) ?
                  (|reg363) : (-reg345)) * $unsigned((reg363 ?
                  reg371 : reg344)))));
              reg375 = (wire311 ?
                  $signed("KnQyfcWn3s") : reg359[(4'h9):(3'h4)]);
              reg376 <= (^($unsigned(($unsigned(reg327) >>> $unsigned((8'hbe)))) > $unsigned((8'hb8))));
            end
          reg377 = (($signed(("" ?
                  (reg337 ?
                      reg373 : reg372) : (~forvar346))) || reg372[(4'hc):(1'h1)]) ?
              (!$unsigned({reg334[(2'h2):(2'h2)],
                  $signed((8'ha3))})) : reg323[(1'h0):(1'h0)]);
          for (forvar378 = (1'h0); (forvar378 < (2'h3)); forvar378 = (forvar378 + (1'h1)))
            begin
              reg379 = (((($signed(reg344) || (reg338 ?
                      reg344 : reg376)) > $signed((~^forvar346))) ?
                  $signed(forvar341[(4'h8):(1'h0)]) : ((~&(reg363 ?
                          reg351 : reg339)) ?
                      wire314[(1'h1):(1'h0)] : $signed((-forvar367)))) == ((+(8'hb2)) ?
                  reg315[(5'h11):(3'h6)] : reg335));
              reg380 <= {$unsigned((^~$unsigned(((7'h43) > reg371))))};
              reg381 = reg351;
              reg382 = (~^forvar341);
            end
          if (({$unsigned({(reg344 >= (8'ha7))}),
              ($signed($signed((7'h43))) ?
                  ((forvar348 ? reg354 : wire309) ?
                      $signed(wire314) : ((8'hb9) != reg330)) : $signed((7'h41)))} >> $unsigned(("xhxsf0P1iQlDRUBz9lH" ?
              (^(^reg363)) : reg352))))
            begin
              reg383 <= {(^(^reg381)), (^$unsigned((~$unsigned(reg334))))};
              reg384 <= $signed(((($unsigned(reg372) ?
                      reg375[(2'h3):(1'h0)] : (-reg330)) >> ($signed(reg352) + forvar353)) ?
                  {reg345[(3'h7):(1'h0)],
                      (!$signed(reg364))} : $unsigned({wire310[(2'h3):(1'h1)],
                      (reg353 ? reg375 : reg364)})));
              reg385 <= (+$unsigned((((reg363 + reg344) >> (reg342 == reg349)) < ($signed((8'had)) ?
                  (reg361 ? forvar378 : forvar341) : reg375[(5'h12):(3'h5)]))));
            end
          else
            begin
              reg383 <= {$unsigned((&(8'ha6)))};
              reg384 <= (8'hbc);
              reg385 <= wire309[(2'h2):(2'h2)];
            end
        end
    end
  assign wire386 = $signed($unsigned((|$unsigned({reg354}))));
  assign wire387 = (8'hbb);
  assign wire388 = {reg385, reg350[(1'h1):(1'h0)]};
  assign wire389 = $signed(reg342);
  always
    @(posedge clk) begin
      if ($signed($signed($signed(wire310))))
        begin
          for (forvar390 = (1'h0); (forvar390 < (1'h0)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 <= ($unsigned(({(&reg358),
                      {(8'ha8)}} * ($unsigned(reg357) ?
                      ((8'hbf) ? reg325 : wire314) : "w"))) ?
                  (reg365[(5'h10):(4'h9)] <<< ($unsigned((reg323 ?
                      reg368 : reg332)) ^ ((reg330 << reg365) <<< $signed((8'haf))))) : (reg334 ?
                      $signed((wire313 ? "RT" : reg323)) : reg324));
              reg392 = reg371;
            end
          reg393 = ({reg319} ?
              reg384[(1'h1):(1'h1)] : $signed($unsigned($signed($unsigned((8'hb7))))));
          reg394 <= (({{{reg348}, ((8'hbb) ? (8'hb6) : reg353)},
              reg352[(4'hb):(1'h0)]} ^ $signed((8'hb5))) >> (8'hb0));
        end
      else
        begin
          for (forvar390 = (1'h0); (forvar390 < (3'h4)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 <= (^reg348);
              reg392 = ((reg323 ?
                  (reg354 >= ($signed(reg385) >= (reg383 * reg339))) : (((^~reg394) && {reg342,
                          reg323}) ?
                      wire314 : $unsigned($unsigned(reg339)))) & wire386[(3'h4):(1'h0)]);
              reg393 = $unsigned(reg374);
              reg394 <= $signed(wire389);
              reg395 <= ($unsigned(($unsigned(reg319) ^~ (reg353 ?
                  (+reg368) : (reg342 ?
                      reg337 : reg332)))) ^ (wire313[(3'h6):(2'h2)] <<< ($signed((reg348 ^~ reg328)) >>> reg357[(3'h7):(2'h3)])));
            end
          reg396 <= (+(8'haf));
        end
      for (forvar397 = (1'h0); (forvar397 < (1'h0)); forvar397 = (forvar397 + (1'h1)))
        begin
          if ((~&reg347))
            begin
              reg398 <= ((("CkcsDL9" ?
                  ($signed(reg360) << (&reg392)) : $unsigned({reg380})) << reg355) || ($unsigned(reg354) ?
                  reg352 : (~|(reg347 ?
                      $signed(wire314) : reg337[(2'h2):(1'h1)]))));
              reg399 = "psWqkDg11B";
              reg400 <= "kEmA1gOINOlgSNxKK";
              reg401 <= {$unsigned(wire389[(3'h4):(3'h4)])};
              reg402 = (^reg376);
            end
          else
            begin
              reg399 = (!$unsigned(($unsigned(reg324[(1'h0):(1'h0)]) ?
                  reg398[(2'h2):(1'h0)] : {$unsigned(reg396)})));
            end
          if ($unsigned(((((~reg399) - reg337[(1'h1):(1'h0)]) <= reg335[(3'h6):(1'h1)]) ?
              reg334 : ($unsigned((-(8'hbc))) ? wire311 : $signed(reg383)))))
            begin
              reg403 <= (~^((~|($unsigned(reg353) == reg354[(1'h0):(1'h0)])) ?
                  (!reg380) : {reg354}));
              reg404 = (~wire312);
              reg405 <= (~^$unsigned((-$unsigned(reg323))));
              reg406 <= $signed(reg337);
              reg407 = (reg328 >= (~wire312));
            end
          else
            begin
              reg403 <= $signed((forvar397 + (~($signed(wire311) ?
                  {reg319} : $unsigned(reg327)))));
            end
          if ((~reg364[(4'hd):(1'h1)]))
            begin
              reg408 = (reg401[(4'ha):(4'ha)] ?
                  reg369 : (forvar390 >> $signed(reg373)));
            end
          else
            begin
              reg408 = reg403;
              reg409 = $unsigned({(|{(reg335 <= reg406), "DUd7"}), "G"});
              reg410 <= (!((~|wire386[(2'h3):(1'h0)]) ?
                  {($unsigned(reg392) ? {reg357, (8'h9d)} : (8'ha5)),
                      $signed({wire311, wire314})} : reg394));
              reg411 <= (8'ha8);
              reg412 = (^($signed(($signed(reg353) >>> (~|reg391))) ?
                  $unsigned(reg339[(1'h1):(1'h0)]) : $signed(($unsigned(reg337) ?
                      $signed((7'h40)) : (reg357 ? reg369 : reg339)))));
            end
          reg413 <= reg368[(4'ha):(1'h1)];
        end
      reg414 <= (((((-reg400) ?
                  (reg342 ? reg353 : (7'h42)) : (|reg358)) >> (7'h42)) ?
              $unsigned(wire309[(4'hb):(3'h4)]) : (wire388 ?
                  ((reg400 && reg332) ?
                      $signed(reg325) : $signed(reg324)) : $unsigned(reg332))) ?
          wire386 : $signed(reg348[(2'h2):(1'h1)]));
    end
  assign wire415 = {$unsigned({(^(reg347 >= reg411)), reg360}),
                       (&$unsigned({(!wire386), reg324[(1'h0):(1'h0)]}))};
  always
    @(posedge clk) begin
      reg416 = (&reg414);
      for (forvar417 = (1'h0); (forvar417 < (1'h1)); forvar417 = (forvar417 + (1'h1)))
        begin
          for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
            begin
              reg419 = wire389;
            end
          reg420 <= {reg394,
              (reg405[(5'h10):(4'hd)] ? $signed((|(^~(8'hb6)))) : reg334)};
          reg421 = $signed($unsigned(("RLnF" ?
              ($unsigned(reg410) - reg319) : $signed((~reg380)))));
        end
      for (forvar422 = (1'h0); (forvar422 < (3'h4)); forvar422 = (forvar422 + (1'h1)))
        begin
          for (forvar423 = (1'h0); (forvar423 < (1'h0)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 = $signed((reg411[(1'h0):(1'h0)] ?
                  ($signed($signed(reg364)) ?
                      ($unsigned((8'ha0)) << (forvar423 ?
                          wire309 : reg368)) : (!"")) : {{{(8'ha2)},
                          (7'h41)}}));
              reg425 = (^~{$unsigned(({(8'hb0)} - $signed(reg330)))});
              reg426 = $signed(reg339);
              reg427 = (7'h43);
              reg428 <= reg335[(3'h5):(1'h1)];
            end
        end
      reg429 = (($unsigned($signed($unsigned(reg391))) && $unsigned(reg398[(4'hd):(3'h4)])) ?
          wire314 : $unsigned(((8'hbd) ?
              $unsigned((wire309 ? reg337 : (8'ha3))) : (+(8'ha7)))));
      for (forvar430 = (1'h0); (forvar430 < (3'h4)); forvar430 = (forvar430 + (1'h1)))
        begin
          reg431 <= ({reg395,
              reg348[(2'h2):(1'h0)]} >> (&(reg358[(3'h6):(3'h5)] >= $unsigned(reg405[(4'h8):(1'h0)]))));
          for (forvar432 = (1'h0); (forvar432 < (1'h0)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= $signed(($unsigned((reg323[(2'h2):(1'h1)] <<< reg405)) >= {(~$signed(wire387))}));
              reg434 = (($unsigned("hXsQKTQ") ?
                      reg337 : reg384[(4'h8):(3'h4)]) ?
                  wire387[(3'h7):(3'h5)] : ((reg332[(3'h5):(2'h3)] >>> (8'hab)) <= wire386[(2'h3):(1'h1)]));
              reg435 <= forvar423[(5'h14):(4'h8)];
              reg436 <= {{$unsigned(((reg413 * reg435) ?
                          $unsigned(reg323) : (reg419 == reg384))),
                      $unsigned($unsigned((wire388 ? reg337 : forvar423)))}};
            end
          reg437 <= reg373;
          for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
            begin
              reg439 = ((forvar418[(4'h9):(4'h9)] || reg383) + reg411[(3'h5):(1'h0)]);
              reg440 <= $unsigned((~|reg380));
              reg441 <= $unsigned(reg398[(1'h0):(1'h0)]);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module103
#(parameter param266 = (({(((8'hb0) >> (8'hb8)) << (~(8'ha1)))} ? (({(8'had), (8'hb0)} ? (^~(8'hb1)) : (8'h9d)) | ({(8'haf)} <= ((8'hb1) ? (8'ha9) : (8'hb6)))) : (((+(8'hab)) ? ((8'haa) ? (8'hb7) : (7'h43)) : ((8'hac) ? (8'had) : (8'h9c))) ? (8'ha0) : (+((8'ha6) ? (8'hbc) : (8'h9f))))) ? ((8'hac) ? ((!((8'hb0) ~^ (8'h9f))) ? {((7'h42) ? (8'hb4) : (8'hbb))} : (((8'hb8) ? (8'ha3) : (8'ha0)) >>> ((8'h9c) ? (8'ha7) : (8'hba)))) : (&(^~((8'ha1) - (8'had))))) : ((~&(((8'ha7) ? (8'hb8) : (8'hb7)) ? {(8'h9f)} : (-(8'ha5)))) ? (~&({(8'ha3)} >>> ((8'hb3) <= (8'ha1)))) : (^~(((8'ha6) ? (8'hb7) : (8'h9e)) | (!(8'ha7)))))))
(y, clk, wire107, wire106, wire105, wire104);
  output wire [(32'h721):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire107;
  input wire [(3'h7):(1'h0)] wire106;
  input wire [(5'h13):(1'h0)] wire105;
  input wire signed [(3'h7):(1'h0)] wire104;
  wire signed [(5'h15):(1'h0)] wire265;
  wire signed [(4'h9):(1'h0)] wire264;
  wire signed [(4'hb):(1'h0)] wire263;
  wire signed [(2'h2):(1'h0)] wire216;
  wire signed [(5'h10):(1'h0)] wire215;
  wire [(5'h14):(1'h0)] wire214;
  wire signed [(4'hc):(1'h0)] wire172;
  wire [(5'h10):(1'h0)] wire136;
  wire [(4'hb):(1'h0)] wire135;
  wire [(5'h14):(1'h0)] wire134;
  wire [(4'hc):(1'h0)] wire133;
  wire signed [(5'h12):(1'h0)] wire120;
  wire signed [(5'h14):(1'h0)] wire108;
  reg signed [(4'hf):(1'h0)] reg262 = (1'h0);
  reg [(5'h14):(1'h0)] reg261 = (1'h0);
  reg [(3'h6):(1'h0)] reg258 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg257 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg252 = (1'h0);
  reg [(2'h3):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg249 = (1'h0);
  reg [(3'h5):(1'h0)] reg247 = (1'h0);
  reg [(4'ha):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg244 = (1'h0);
  reg [(4'he):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg242 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg240 = (1'h0);
  reg [(5'h15):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg [(4'hc):(1'h0)] reg236 = (1'h0);
  reg [(4'hf):(1'h0)] reg235 = (1'h0);
  reg [(4'hd):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg226 = (1'h0);
  reg [(5'h11):(1'h0)] reg224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg222 = (1'h0);
  reg signed [(4'he):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg210 = (1'h0);
  reg [(4'hc):(1'h0)] reg209 = (1'h0);
  reg [(2'h3):(1'h0)] reg207 = (1'h0);
  reg [(5'h15):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg204 = (1'h0);
  reg [(4'hd):(1'h0)] reg201 = (1'h0);
  reg [(5'h11):(1'h0)] reg200 = (1'h0);
  reg [(4'h9):(1'h0)] reg195 = (1'h0);
  reg [(5'h13):(1'h0)] reg194 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg193 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg188 = (1'h0);
  reg [(5'h15):(1'h0)] reg187 = (1'h0);
  reg [(4'h8):(1'h0)] reg182 = (1'h0);
  reg [(3'h4):(1'h0)] reg180 = (1'h0);
  reg [(3'h5):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg177 = (1'h0);
  reg [(3'h6):(1'h0)] reg174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg171 = (1'h0);
  reg [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg164 = (1'h0);
  reg [(5'h15):(1'h0)] reg163 = (1'h0);
  reg [(5'h15):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg154 = (1'h0);
  reg [(4'hc):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg151 = (1'h0);
  reg [(3'h5):(1'h0)] reg140 = (1'h0);
  reg [(4'hb):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg132 = (1'h0);
  reg [(5'h12):(1'h0)] reg128 = (1'h0);
  reg [(4'he):(1'h0)] reg126 = (1'h0);
  reg signed [(4'he):(1'h0)] reg122 = (1'h0);
  reg [(5'h14):(1'h0)] reg121 = (1'h0);
  reg [(4'hf):(1'h0)] reg118 = (1'h0);
  reg [(4'hb):(1'h0)] reg116 = (1'h0);
  reg [(2'h2):(1'h0)] reg114 = (1'h0);
  reg [(5'h13):(1'h0)] reg113 = (1'h0);
  reg [(4'hb):(1'h0)] reg110 = (1'h0);
  reg [(3'h6):(1'h0)] reg260 = (1'h0);
  reg [(2'h3):(1'h0)] reg259 = (1'h0);
  reg [(4'hf):(1'h0)] reg256 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg254 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar251 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg246 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar241 = (1'h0);
  reg [(5'h11):(1'h0)] forvar239 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar234 = (1'h0);
  reg [(4'h9):(1'h0)] reg231 = (1'h0);
  reg [(3'h7):(1'h0)] reg230 = (1'h0);
  reg [(3'h5):(1'h0)] forvar229 = (1'h0);
  reg [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'hc):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg220 = (1'h0);
  reg [(3'h6):(1'h0)] forvar219 = (1'h0);
  reg [(4'hd):(1'h0)] reg218 = (1'h0);
  reg [(3'h4):(1'h0)] reg213 = (1'h0);
  reg [(5'h12):(1'h0)] reg212 = (1'h0);
  reg [(4'ha):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar208 = (1'h0);
  reg [(4'hc):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar202 = (1'h0);
  reg [(4'h8):(1'h0)] forvar199 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg197 = (1'h0);
  reg [(5'h10):(1'h0)] forvar196 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar193 = (1'h0);
  reg [(3'h7):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg190 = (1'h0);
  reg [(4'ha):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg186 = (1'h0);
  reg [(2'h2):(1'h0)] reg185 = (1'h0);
  reg [(2'h2):(1'h0)] reg184 = (1'h0);
  reg [(4'he):(1'h0)] forvar183 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg181 = (1'h0);
  reg [(4'hd):(1'h0)] reg179 = (1'h0);
  reg [(4'he):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar175 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg173 = (1'h0);
  reg [(5'h14):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg168 = (1'h0);
  reg [(3'h7):(1'h0)] forvar166 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg165 = (1'h0);
  reg [(5'h11):(1'h0)] reg162 = (1'h0);
  reg [(4'hf):(1'h0)] reg160 = (1'h0);
  reg [(4'hd):(1'h0)] forvar159 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar158 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg157 = (1'h0);
  reg [(2'h3):(1'h0)] reg156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg152 = (1'h0);
  reg [(4'hf):(1'h0)] forvar150 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg149 = (1'h0);
  reg [(5'h12):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg144 = (1'h0);
  reg [(2'h2):(1'h0)] forvar143 = (1'h0);
  reg [(5'h11):(1'h0)] reg142 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg141 = (1'h0);
  reg [(4'h8):(1'h0)] reg138 = (1'h0);
  reg [(4'hb):(1'h0)] forvar137 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg131 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg130 = (1'h0);
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  reg [(4'ha):(1'h0)] reg127 = (1'h0);
  reg [(3'h4):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar124 = (1'h0);
  reg [(4'h8):(1'h0)] forvar123 = (1'h0);
  reg [(3'h6):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar117 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg115 = (1'h0);
  reg [(4'h8):(1'h0)] forvar112 = (1'h0);
  reg [(5'h12):(1'h0)] forvar111 = (1'h0);
  reg [(4'h8):(1'h0)] reg109 = (1'h0);
  assign y = {wire265,
                 wire264,
                 wire263,
                 wire216,
                 wire215,
                 wire214,
                 wire172,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire120,
                 wire108,
                 reg262,
                 reg261,
                 reg258,
                 reg257,
                 reg253,
                 reg252,
                 reg250,
                 reg249,
                 reg247,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg240,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg233,
                 reg232,
                 reg226,
                 reg224,
                 reg222,
                 reg221,
                 reg217,
                 reg210,
                 reg209,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg201,
                 reg200,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg188,
                 reg187,
                 reg182,
                 reg180,
                 reg178,
                 reg177,
                 reg174,
                 reg171,
                 reg169,
                 reg167,
                 reg164,
                 reg163,
                 reg161,
                 reg155,
                 reg154,
                 reg153,
                 reg151,
                 reg140,
                 reg139,
                 reg137,
                 reg132,
                 reg128,
                 reg126,
                 reg122,
                 reg121,
                 reg118,
                 reg116,
                 reg114,
                 reg113,
                 reg110,
                 reg260,
                 reg259,
                 reg256,
                 reg255,
                 reg254,
                 forvar251,
                 reg248,
                 reg246,
                 forvar241,
                 forvar239,
                 forvar234,
                 reg231,
                 reg230,
                 forvar229,
                 reg228,
                 reg227,
                 reg225,
                 reg223,
                 reg220,
                 forvar219,
                 reg218,
                 reg213,
                 reg212,
                 reg211,
                 forvar208,
                 reg203,
                 forvar202,
                 forvar199,
                 reg198,
                 reg197,
                 forvar196,
                 forvar193,
                 reg191,
                 reg190,
                 reg189,
                 reg186,
                 reg185,
                 reg184,
                 forvar183,
                 reg181,
                 reg179,
                 reg176,
                 forvar175,
                 reg173,
                 reg170,
                 reg168,
                 forvar166,
                 reg165,
                 reg162,
                 reg160,
                 forvar159,
                 forvar158,
                 reg157,
                 reg156,
                 reg152,
                 forvar150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 reg141,
                 reg138,
                 forvar137,
                 reg131,
                 reg130,
                 reg129,
                 reg127,
                 reg125,
                 forvar124,
                 forvar123,
                 reg119,
                 forvar117,
                 reg115,
                 forvar112,
                 forvar111,
                 reg109,
                 (1'h0)};
  assign wire108 = (~&$signed((((-wire104) != (|wire104)) && $unsigned(((8'ha3) ?
                       wire107 : wire106)))));
  always
    @(posedge clk) begin
      reg109 = wire106;
      reg110 <= "plgVuTik0D0rLeh";
      for (forvar111 = (1'h0); (forvar111 < (1'h0)); forvar111 = (forvar111 + (1'h1)))
        begin
          for (forvar112 = (1'h0); (forvar112 < (2'h2)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= (~|($unsigned(((wire105 ? forvar111 : (8'haa)) ?
                      (^~forvar111) : wire106[(3'h7):(2'h3)])) ?
                  wire107 : ($unsigned($signed(wire106)) >> forvar112)));
            end
          if ({wire107[(4'h8):(3'h5)]})
            begin
              reg114 <= reg113;
            end
          else
            begin
              reg115 = {(reg110 ?
                      ({(^reg109)} ?
                          (^~{wire106,
                              wire108}) : $unsigned((wire106 != reg110))) : $unsigned((!(reg109 ?
                          reg109 : reg110))))};
              reg116 <= (("fW" ?
                      wire105 : {((forvar112 & wire108) == "IUkrkDfYLqImoYE"),
                          wire106}) ?
                  (8'hb4) : forvar111);
            end
          for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= ($unsigned(wire108) ?
                  wire105[(5'h12):(4'hd)] : (!$unsigned((-$signed(reg116)))));
            end
          reg119 = ({(~^((wire104 ~^ wire108) >> $unsigned(forvar112))),
              $unsigned("h")} && $signed("TmHJSN"));
        end
    end
  assign wire120 = reg118;
  always
    @(posedge clk) begin
      reg121 <= {(~|(^~(~(^~reg116)))), reg118[(2'h2):(1'h0)]};
      reg122 <= ({((-{(8'hbe)}) ? $signed((~&reg114)) : $unsigned((&reg114))),
              ((~|(wire106 ? (7'h41) : reg113)) ?
                  wire120[(4'hc):(4'ha)] : reg118[(3'h6):(2'h3)])} ?
          $signed($unsigned($signed((reg110 * wire108)))) : (reg114 ?
              (~$signed($unsigned((7'h40)))) : (wire108 | {{(8'hb0), wire105},
                  $signed(reg116)})));
      for (forvar123 = (1'h0); (forvar123 < (3'h4)); forvar123 = (forvar123 + (1'h1)))
        begin
          for (forvar124 = (1'h0); (forvar124 < (2'h3)); forvar124 = (forvar124 + (1'h1)))
            begin
              reg125 = ($signed($signed(wire104[(3'h4):(2'h3)])) ?
                  wire107 : ((reg110[(4'ha):(3'h7)] > (~&reg113[(3'h7):(3'h7)])) ?
                      forvar123 : (reg118 ?
                          reg116 : ($unsigned(wire120) - (wire108 && reg113)))));
            end
          if (wire120)
            begin
              reg126 <= (((~&"GI7sRbcH") ?
                      reg121 : ({(forvar124 | reg114)} ?
                          $unsigned(reg122) : reg125)) ?
                  ((((~wire106) ?
                      (-reg122) : $unsigned(forvar124)) * forvar123[(3'h5):(2'h3)]) != $unsigned(((~|(8'haf)) >>> $signed(forvar123)))) : $signed((-forvar124)));
            end
          else
            begin
              reg127 = ((((+$signed(wire104)) ?
                      (~&$signed((7'h44))) : reg110[(3'h7):(2'h2)]) ?
                  ($unsigned((wire107 == wire108)) ?
                      $unsigned("o20dnolBd") : {((7'h44) ~^ reg122),
                          (wire107 + wire108)}) : $unsigned(($signed(reg121) ?
                      $unsigned((8'hbd)) : $unsigned((8'h9d))))) || reg110);
              reg128 <= wire120[(4'hf):(1'h1)];
              reg129 = (wire120 ? reg118[(3'h4):(2'h3)] : reg114);
              reg130 = $unsigned((($unsigned((wire120 == forvar124)) ?
                      (-(reg128 ? wire120 : wire106)) : ($unsigned(reg122) ?
                          $signed(reg122) : (wire104 ? reg114 : reg125))) ?
                  (({reg110} < $unsigned(wire120)) ?
                      reg116[(4'hb):(4'hb)] : (((8'ha3) >= (8'hbd)) ^ ((8'h9e) && reg127))) : "Mu94NTdvXF"));
              reg131 = (~^(wire120 + (wire120[(5'h10):(4'hf)] * ($signed(reg110) << (reg122 ?
                  reg125 : wire104)))));
            end
          reg132 <= (((wire104[(1'h1):(1'h0)] >= ({reg125} ~^ (&forvar124))) || ((!(reg131 ?
              reg113 : reg129)) != (!(reg122 ^~ (8'hba))))) >= (-wire106[(3'h4):(1'h1)]));
        end
    end
  assign wire133 = ((((((7'h41) ? reg116 : (8'hba)) ?
                           (reg118 >> wire120) : $unsigned((8'hb5))) ?
                       ((reg128 ? reg128 : wire104) ?
                           (reg113 <<< reg113) : reg118) : $unsigned((reg132 ^~ (8'hb4)))) + reg121) != reg110[(4'ha):(4'h9)]);
  assign wire134 = {wire105, reg121};
  assign wire135 = {{$unsigned(("yyJQOYJWQTUm3Rb8cvnX" ?
                               $unsigned(wire133) : (~&wire104)))},
                       reg126[(4'hc):(1'h1)]};
  assign wire136 = $signed(reg116);
  always
    @(posedge clk) begin
      if (wire135[(1'h1):(1'h1)])
        begin
          for (forvar137 = (1'h0); (forvar137 < (2'h2)); forvar137 = (forvar137 + (1'h1)))
            begin
              reg138 = "gO0W3RTif";
            end
        end
      else
        begin
          if ($unsigned($unsigned(wire104[(2'h3):(2'h2)])))
            begin
              reg137 <= {(&"alF2DSsiCT")};
              reg138 = $signed(wire104[(3'h6):(1'h0)]);
              reg139 <= $unsigned((|wire105[(5'h11):(3'h6)]));
              reg140 <= (7'h44);
            end
          else
            begin
              reg137 <= wire136;
              reg139 <= (8'hb7);
              reg140 <= wire136[(4'hf):(4'ha)];
              reg141 = {{reg118, forvar137}};
              reg142 = reg128[(4'hf):(3'h6)];
            end
          for (forvar143 = (1'h0); (forvar143 < (1'h1)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 = reg137[(2'h3):(1'h0)];
              reg145 = reg144;
              reg146 = $unsigned($unsigned((wire120 ?
                  $unsigned("sLOxBt10iP1KrW3BS2L") : ({(8'hb5),
                      reg113} != reg121))));
              reg147 = $signed(reg145[(2'h3):(2'h3)]);
              reg148 = $unsigned($signed(($unsigned({reg121,
                  wire108}) ^ (!(-reg137)))));
            end
          reg149 = $unsigned(reg114);
        end
      for (forvar150 = (1'h0); (forvar150 < (2'h3)); forvar150 = (forvar150 + (1'h1)))
        begin
          if (($unsigned((~&reg147[(2'h2):(2'h2)])) ^~ {wire105,
              reg128[(4'hf):(2'h2)]}))
            begin
              reg151 <= (8'ha4);
              reg152 = reg146[(2'h3):(1'h0)];
            end
          else
            begin
              reg151 <= "kSWZvhw";
              reg153 <= reg110;
              reg154 <= wire134;
              reg155 <= (~^$signed((reg154 ?
                  $unsigned((reg154 <= reg147)) : {(~reg144),
                      reg137[(4'hf):(4'h8)]})));
            end
          reg156 = reg138[(2'h3):(2'h3)];
        end
      reg157 = ((((^~reg144[(3'h6):(2'h3)]) > $unsigned((wire105 ?
              (7'h40) : wire107))) == $unsigned(wire104[(3'h7):(3'h4)])) ?
          reg113[(4'h9):(2'h3)] : {({((8'ha6) < (8'ha8)),
                  $unsigned(reg147)} + ((reg154 ? reg110 : wire108) ^ (reg141 ?
                  wire134 : reg141)))});
      for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
        begin
          for (forvar159 = (1'h0); (forvar159 < (3'h4)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 = $unsigned(reg145);
              reg161 <= (!(-(7'h44)));
              reg162 = (-{(!{$signed(reg113), reg154[(2'h2):(2'h2)]}),
                  (8'hbe)});
            end
          if ((reg156 ?
              $unsigned(reg126[(4'h8):(4'h8)]) : {(~$unsigned($signed(reg148)))}))
            begin
              reg163 <= ((reg153 && (($unsigned(wire104) * wire134) > $signed((|reg128)))) || ((~$signed($unsigned(reg152))) ?
                  reg161[(3'h5):(3'h5)] : ($signed(reg118[(4'hc):(4'h9)]) ?
                      $signed($unsigned(wire120)) : reg139[(2'h2):(1'h0)])));
              reg164 <= ({$signed($unsigned((forvar158 ?
                      reg156 : reg163)))} != $unsigned($signed(forvar158)));
              reg165 = $signed((((!$unsigned(reg157)) ?
                      (!"qzoKpAX5X89f") : reg154) ?
                  forvar143[(1'h0):(1'h0)] : reg151[(2'h3):(1'h0)]));
            end
          else
            begin
              reg163 <= $unsigned((8'hb3));
            end
          for (forvar166 = (1'h0); (forvar166 < (1'h1)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= $signed({(8'hbd)});
              reg168 = ((+reg162) * {reg161[(3'h7):(2'h2)]});
              reg169 <= (8'ha1);
              reg170 = reg121;
              reg171 <= (^(|{(reg128 ? (wire135 | reg149) : {reg156})}));
            end
        end
    end
  assign wire172 = ((&(~reg116)) - (({(reg114 ? wire107 : wire106),
                           ((8'haf) >= reg128)} ?
                       ($signed(reg132) > (reg164 ?
                           reg118 : wire136)) : {wire105,
                           reg113[(3'h6):(3'h4)]}) + $unsigned((wire104 ?
                       wire108 : reg151))));
  always
    @(posedge clk) begin
      reg173 = $signed((({$signed((8'hab))} ? wire133 : $signed(reg151)) ?
          reg155 : wire135[(2'h3):(2'h3)]));
      reg174 <= $signed(wire133);
      for (forvar175 = (1'h0); (forvar175 < (1'h1)); forvar175 = (forvar175 + (1'h1)))
        begin
          reg176 = $unsigned({{$signed((7'h44)),
                  $signed((reg167 ? reg110 : reg118))}});
          if ($signed(((~$unsigned({wire105})) ?
              ($signed(reg164[(4'ha):(3'h7)]) ^ (|reg140[(3'h5):(2'h3)])) : wire108)))
            begin
              reg177 <= reg174[(3'h5):(3'h4)];
              reg178 <= $signed(wire107[(3'h6):(3'h5)]);
              reg179 = reg114;
              reg180 <= (("uOwPxv9JUhwWNfLrE6tq" || $signed((+(reg128 ?
                      (7'h42) : (8'ha4))))) ?
                  (({(reg161 ? reg153 : reg174),
                      {wire120}} | {(wire134 >>> reg171)}) ~^ (($unsigned(forvar175) ?
                      (~&wire136) : $unsigned(reg140)) - $unsigned($unsigned(reg128)))) : reg122[(3'h7):(1'h1)]);
              reg181 = reg173;
            end
          else
            begin
              reg179 = (reg121[(5'h10):(4'h9)] ?
                  reg118 : reg177[(2'h3):(2'h2)]);
              reg180 <= (wire106[(1'h1):(1'h1)] || (-wire108[(4'hb):(4'ha)]));
            end
          reg182 <= wire172[(4'ha):(1'h1)];
        end
      for (forvar183 = (1'h0); (forvar183 < (2'h3)); forvar183 = (forvar183 + (1'h1)))
        begin
          if ($signed(wire133))
            begin
              reg184 = $signed(($signed($unsigned((reg140 < reg116))) ?
                  reg126[(3'h6):(1'h0)] : reg169));
              reg185 = {$unsigned(($unsigned($unsigned(reg181)) <<< ""))};
              reg186 = reg185[(2'h2):(2'h2)];
            end
          else
            begin
              reg187 <= $unsigned(((($unsigned((8'ha9)) != reg151) ?
                  $unsigned(wire106) : (^~(^~(8'hb7)))) || $signed(reg154[(1'h1):(1'h1)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg188 <= $unsigned($unsigned((~&wire120[(3'h4):(2'h3)])));
      reg189 = reg154[(1'h1):(1'h1)];
      if (((~&$signed(reg126)) || {(($unsigned(wire134) ?
                  (reg188 ? (8'hb5) : reg189) : reg126[(3'h5):(1'h0)]) ?
              reg154[(3'h5):(3'h4)] : reg128),
          (reg180 ?
              reg116 : (((8'ha0) ? wire136 : wire135) ?
                  (reg137 ? wire106 : reg155) : $unsigned((8'ha9))))}))
        begin
          reg190 = $unsigned($unsigned((8'hac)));
          reg191 = reg122[(2'h3):(1'h1)];
          reg192 <= $unsigned((wire134[(5'h12):(4'ha)] >= reg189[(3'h5):(1'h1)]));
          reg193 <= ($unsigned((reg190[(2'h2):(1'h0)] <= $unsigned(wire133[(2'h3):(2'h3)]))) ?
              reg167[(1'h0):(1'h0)] : ($unsigned($unsigned(reg167)) >= (8'hb5)));
        end
      else
        begin
          reg192 <= (reg113[(5'h12):(4'ha)] != $unsigned(reg128[(1'h1):(1'h0)]));
          for (forvar193 = (1'h0); (forvar193 < (2'h3)); forvar193 = (forvar193 + (1'h1)))
            begin
              reg194 <= reg180;
              reg195 <= (wire107[(1'h0):(1'h0)] ?
                  $unsigned(({"HE5UJM1vT9a3S"} ?
                      (+$signed((8'hbc))) : $signed(reg126))) : $unsigned((wire105[(3'h7):(3'h4)] ?
                      (+reg137[(5'h11):(3'h6)]) : {$unsigned(forvar193)})));
            end
          for (forvar196 = (1'h0); (forvar196 < (3'h4)); forvar196 = (forvar196 + (1'h1)))
            begin
              reg197 = ((~reg195) ? wire172 : forvar196);
              reg198 = (~^(&"GTIuQO3"));
            end
        end
      for (forvar199 = (1'h0); (forvar199 < (1'h1)); forvar199 = (forvar199 + (1'h1)))
        begin
          reg200 <= wire133;
          reg201 <= (8'h9f);
          for (forvar202 = (1'h0); (forvar202 < (1'h1)); forvar202 = (forvar202 + (1'h1)))
            begin
              reg203 = wire134[(2'h3):(2'h3)];
              reg204 <= ($signed((^(reg200 >> (reg192 << (8'hab))))) | $signed((8'hb9)));
              reg205 <= {$signed($unsigned(reg137[(3'h5):(1'h0)])),
                  reg174[(3'h4):(1'h1)]};
              reg206 <= ((8'hb7) ?
                  ({reg205[(2'h3):(1'h1)]} ?
                      (&reg200[(4'hc):(3'h5)]) : (({forvar199} ?
                          (~(8'h9f)) : ((8'h9d) & reg118)) ~^ reg114)) : $signed(reg187));
            end
          reg207 <= ({(wire134 ?
                      $unsigned(forvar193) : ($signed(wire107) ?
                          (reg188 & reg182) : (wire120 == reg140))),
                  ((^~$signed(reg110)) ?
                      reg126[(1'h1):(1'h1)] : (((8'hb6) ?
                          reg163 : wire135) | $signed((8'haf))))} ?
              {(7'h43)} : reg182[(2'h3):(1'h1)]);
          for (forvar208 = (1'h0); (forvar208 < (1'h1)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 <= $unsigned(($unsigned(($signed((8'hb3)) << $unsigned(wire106))) ?
                  ((7'h43) ?
                      (!$unsigned(reg207)) : "eFMniSdb2") : (reg121[(4'he):(4'h9)] | wire106[(3'h7):(3'h4)])));
              reg210 <= reg182;
              reg211 = $unsigned((~^$signed((^$signed(reg118)))));
              reg212 = ((&(8'had)) ?
                  reg153 : {((8'hbb) && forvar199[(2'h3):(2'h3)])});
              reg213 = reg137[(3'h6):(3'h6)];
            end
        end
    end
  assign wire214 = ((|({(~|reg113)} && (8'ha7))) || {reg163[(3'h7):(2'h3)],
                       (&$unsigned($signed((8'ha9))))});
  assign wire215 = $unsigned($unsigned($signed({$unsigned(reg171)})));
  assign wire216 = (+$signed((8'hb6)));
  always
    @(posedge clk) begin
      reg217 <= (&((({wire133} <<< (reg195 <= wire120)) << $signed($unsigned(reg137))) * wire216));
    end
  always
    @(posedge clk) begin
      reg218 = $signed($signed($signed(reg210[(5'h10):(1'h1)])));
    end
  always
    @(posedge clk) begin
      for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
        begin
          if ($signed((^reg155)))
            begin
              reg220 = (reg200 ?
                  reg161 : ($signed(($unsigned(reg171) || (~reg137))) ?
                      (~^(reg182 >= reg210[(3'h7):(1'h0)])) : "zU"));
              reg221 <= reg139[(3'h4):(1'h1)];
              reg222 <= wire106;
            end
          else
            begin
              reg221 <= (!wire104[(3'h7):(1'h1)]);
              reg223 = $unsigned($signed($unsigned($signed((reg121 ?
                  reg201 : reg188)))));
              reg224 <= ("GqkphcizQ" | {$signed({forvar219, wire105}),
                  ({$unsigned(wire106), (wire106 ? (8'hba) : reg194)} ?
                      ($signed((8'h9d)) <= reg167[(1'h1):(1'h0)]) : $signed($signed(reg161)))});
              reg225 = (8'hb7);
              reg226 <= {$signed((-{(~|reg171)}))};
            end
        end
      reg227 = ($signed(reg163) ?
          (~|(wire134 ~^ (~^{(8'h9f),
              reg205}))) : {$signed(reg114[(1'h1):(1'h0)]),
              ((reg174[(3'h4):(2'h2)] < $unsigned((8'hbc))) ?
                  ($signed(reg178) ?
                      ((8'ha9) < (8'ha2)) : $signed(reg195)) : reg201)});
      reg228 = (-$signed(((8'haf) ? $unsigned((-reg223)) : reg192)));
      for (forvar229 = (1'h0); (forvar229 < (3'h4)); forvar229 = (forvar229 + (1'h1)))
        begin
          if ($unsigned($unsigned(reg154)))
            begin
              reg230 = (~&$signed((reg177 ?
                  ($unsigned(reg169) ?
                      {reg118, wire134} : reg180) : (|reg122))));
              reg231 = (!($unsigned((^(|reg114))) ?
                  {$unsigned(reg174)} : reg187));
            end
          else
            begin
              reg232 <= "bp1dL2RqpMy";
              reg233 <= (~&(({$unsigned(reg193)} >>> (-(wire135 ^ (8'ha4)))) >= ((~(reg195 <= reg187)) ?
                  {$unsigned(reg154),
                      "GsRHE3PagDQxKw7K8U"} : (|(reg140 >= reg222)))));
            end
          for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= ($unsigned(($unsigned(reg140) ?
                      $signed((~reg232)) : $unsigned("CQC86K992VEdumA"))) ?
                  $signed(reg169[(3'h6):(2'h2)]) : (8'ha7));
            end
          reg236 <= reg140[(3'h5):(3'h5)];
          reg237 <= $unsigned((reg132 ?
              forvar219[(3'h5):(1'h0)] : ($signed($signed((8'ha8))) ?
                  (reg205 >>> reg139[(4'hb):(1'h0)]) : (8'hbd))));
        end
    end
  always
    @(posedge clk) begin
      reg238 <= ($signed(reg177[(3'h5):(3'h5)]) << $unsigned((wire120[(1'h0):(1'h0)] ?
          reg151[(2'h3):(2'h3)] : reg137[(2'h2):(2'h2)])));
      for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
        begin
          reg240 <= reg194;
          for (forvar241 = (1'h0); (forvar241 < (3'h4)); forvar241 = (forvar241 + (1'h1)))
            begin
              reg242 <= ({((8'ha9) || forvar239[(4'hd):(4'h8)])} && (8'ha1));
              reg243 <= (~&$signed({$unsigned((reg192 | reg200))}));
              reg244 <= {reg192[(1'h1):(1'h0)], reg209[(2'h2):(2'h2)]};
              reg245 <= ($unsigned((~^reg224)) ?
                  (((-(reg137 >= reg155)) & (&$unsigned(reg205))) ?
                      ({wire172[(3'h4):(2'h2)]} ?
                          ((wire107 ^~ (8'haa)) | (reg221 ?
                              wire136 : (8'hbc))) : ($unsigned((8'hbf)) <= $signed(wire136))) : ($unsigned($unsigned(reg164)) ?
                          {$signed((8'hab)),
                              $signed(reg132)} : {reg238[(4'h9):(1'h1)],
                              reg137})) : $signed((^($unsigned(reg240) <= reg187[(3'h4):(2'h3)]))));
            end
          if ((((8'hb4) ^ $signed((8'hb6))) ^~ (7'h42)))
            begin
              reg246 = {{((-$signed(reg140)) ?
                          $unsigned({reg232}) : $unsigned(reg174)),
                      $unsigned((~&(|reg161)))}};
            end
          else
            begin
              reg247 <= reg193;
              reg248 = ($signed(($signed(reg222) & (-reg163[(5'h15):(4'hd)]))) ?
                  $signed(reg247[(1'h1):(1'h1)]) : reg182);
              reg249 <= reg126[(4'hc):(4'h9)];
            end
          reg250 <= (($signed(((wire135 ~^ reg114) ?
              wire172[(2'h3):(1'h1)] : wire120)) >>> (&reg221)) >= ((^$signed(reg210[(5'h13):(5'h11)])) < $signed((~|$signed(reg174)))));
        end
      for (forvar251 = (1'h0); (forvar251 < (2'h3)); forvar251 = (forvar251 + (1'h1)))
        begin
          if ($signed(forvar251[(1'h0):(1'h0)]))
            begin
              reg252 <= reg195;
              reg253 <= {(8'hbd)};
            end
          else
            begin
              reg254 = ($unsigned(wire136[(4'hd):(3'h7)]) ?
                  $signed(reg245) : $signed(($signed($signed((8'haf))) >>> {wire214})));
              reg255 = ((~{((~^reg167) ? reg116 : reg243[(4'ha):(2'h2)]),
                  (|(^wire215))}) != ((((reg151 << reg169) >= $unsigned(reg238)) - reg206) ?
                  (((reg114 ?
                      (8'haf) : wire214) | (reg163 != reg222)) <= "CPEx") : ((|reg236[(1'h1):(1'h1)]) ?
                      "rVdkm4ktcD" : ((reg245 >>> (8'ha9)) ?
                          wire134 : (^~wire214)))));
              reg256 = ((~|$signed($unsigned((&reg222)))) ~^ $unsigned($signed(reg243)));
              reg257 <= ((^~{({reg180, reg153} ? $signed(reg217) : reg116),
                      (^~reg163)}) ?
                  (($signed((reg171 | reg209)) - ((reg232 + wire136) ?
                          {(8'haf)} : ((8'hab) ? reg153 : reg255))) ?
                      (reg161 ^~ ({reg233} | reg254[(3'h6):(1'h1)])) : ((~&(&reg161)) ?
                          $unsigned((|(8'haa))) : (~^((8'hb8) == reg210)))) : $unsigned(reg180));
              reg258 <= {"TkJzUBemmbwNQzpSr"};
            end
          reg259 = (reg118 >= reg180);
          reg260 = (^(~&$signed($unsigned($unsigned(reg194)))));
          reg261 <= $signed(reg122);
        end
      reg262 <= $signed((~^(reg177[(1'h1):(1'h1)] << (~$signed(reg118)))));
    end
  assign wire263 = reg209;
  assign wire264 = {(~|{reg161}), {wire135}};
  assign wire265 = (reg171 ?
                       (+reg224[(4'hf):(2'h2)]) : ($signed((((8'hb1) ^ reg249) ?
                               reg201[(3'h6):(3'h5)] : reg240[(2'h2):(2'h2)])) ?
                           wire104 : ($unsigned((reg237 ? reg233 : (8'hb7))) ?
                               ((^reg244) ?
                                   reg247[(3'h4):(2'h3)] : wire214) : wire120)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module19
#(parameter param99 = (({(((7'h40) ? (7'h43) : (7'h43)) == {(8'hb9)})} & ((~(|(8'hb6))) ? (|(~&(8'ha2))) : (((8'haf) ^~ (8'ha2)) ? {(8'had)} : {(8'ha8)}))) < (({(-(8'hba))} ? {{(8'hb7)}, ((8'hbf) ? (8'hba) : (8'hbe))} : {(~(7'h42))}) | ((~&((8'hae) ? (8'hb2) : (8'h9c))) ? (~^((8'ha8) ? (8'ha4) : (8'h9f))) : (~|(~^(8'hbf)))))), 
parameter param100 = (param99 & ((|({param99} < param99)) ? (((param99 ? param99 : param99) >> param99) ? (~^(8'hbc)) : {((8'hb0) ? param99 : param99), ((8'hb6) ? (7'h44) : param99)}) : (^~(8'ha7)))))
(y, clk, wire23, wire22, wire21, wire20);
  output wire [(32'h34d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire23;
  input wire signed [(5'h11):(1'h0)] wire22;
  input wire signed [(4'hd):(1'h0)] wire21;
  input wire signed [(5'h15):(1'h0)] wire20;
  wire signed [(5'h14):(1'h0)] wire71;
  wire signed [(3'h4):(1'h0)] wire70;
  wire signed [(3'h4):(1'h0)] wire61;
  wire signed [(5'h11):(1'h0)] wire60;
  wire [(4'hd):(1'h0)] wire37;
  wire [(4'hd):(1'h0)] wire26;
  wire [(4'h8):(1'h0)] wire24;
  reg signed [(5'h10):(1'h0)] reg97 = (1'h0);
  reg signed [(4'he):(1'h0)] reg94 = (1'h0);
  reg [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg91 = (1'h0);
  reg [(4'h9):(1'h0)] reg89 = (1'h0);
  reg [(4'h9):(1'h0)] reg87 = (1'h0);
  reg [(4'ha):(1'h0)] reg85 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg80 = (1'h0);
  reg [(4'ha):(1'h0)] reg79 = (1'h0);
  reg [(4'h8):(1'h0)] reg76 = (1'h0);
  reg [(5'h13):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg67 = (1'h0);
  reg [(5'h13):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg64 = (1'h0);
  reg [(3'h4):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg57 = (1'h0);
  reg [(4'he):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg51 = (1'h0);
  reg [(4'hd):(1'h0)] reg49 = (1'h0);
  reg [(4'hb):(1'h0)] reg48 = (1'h0);
  reg [(3'h6):(1'h0)] reg47 = (1'h0);
  reg [(3'h4):(1'h0)] reg45 = (1'h0);
  reg [(4'hc):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg27 = (1'h0);
  reg [(4'hc):(1'h0)] reg25 = (1'h0);
  reg [(5'h10):(1'h0)] reg86 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg98 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg95 = (1'h0);
  reg [(3'h4):(1'h0)] reg93 = (1'h0);
  reg [(2'h2):(1'h0)] reg90 = (1'h0);
  reg [(3'h7):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar86 = (1'h0);
  reg [(2'h2):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar83 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar81 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg78 = (1'h0);
  reg [(5'h13):(1'h0)] reg77 = (1'h0);
  reg [(3'h4):(1'h0)] forvar75 = (1'h0);
  reg [(2'h2):(1'h0)] forvar73 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg69 = (1'h0);
  reg [(4'he):(1'h0)] reg66 = (1'h0);
  reg [(4'hc):(1'h0)] forvar63 = (1'h0);
  reg [(2'h2):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg58 = (1'h0);
  reg [(3'h5):(1'h0)] reg56 = (1'h0);
  reg [(5'h10):(1'h0)] forvar54 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg53 = (1'h0);
  reg [(5'h14):(1'h0)] forvar52 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar50 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar44 = (1'h0);
  reg [(3'h7):(1'h0)] forvar43 = (1'h0);
  reg [(4'h8):(1'h0)] reg42 = (1'h0);
  reg [(5'h13):(1'h0)] reg40 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar39 = (1'h0);
  reg [(5'h13):(1'h0)] forvar38 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg36 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg32 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar31 = (1'h0);
  reg [(5'h12):(1'h0)] reg30 = (1'h0);
  reg [(4'hc):(1'h0)] forvar29 = (1'h0);
  reg [(3'h7):(1'h0)] forvar28 = (1'h0);
  assign y = {wire71,
                 wire70,
                 wire61,
                 wire60,
                 wire37,
                 wire26,
                 wire24,
                 reg97,
                 reg94,
                 reg92,
                 reg91,
                 reg89,
                 reg87,
                 reg85,
                 reg82,
                 reg80,
                 reg79,
                 reg76,
                 reg74,
                 reg68,
                 reg67,
                 reg65,
                 reg64,
                 reg62,
                 reg59,
                 reg57,
                 reg55,
                 reg51,
                 reg49,
                 reg48,
                 reg47,
                 reg45,
                 reg41,
                 reg33,
                 reg27,
                 reg25,
                 reg86,
                 reg98,
                 reg96,
                 reg95,
                 reg93,
                 reg90,
                 reg88,
                 forvar86,
                 reg84,
                 forvar83,
                 forvar81,
                 reg78,
                 reg77,
                 forvar75,
                 forvar73,
                 reg72,
                 reg69,
                 reg66,
                 forvar63,
                 reg63,
                 reg58,
                 reg56,
                 forvar54,
                 reg53,
                 forvar52,
                 forvar50,
                 reg46,
                 forvar44,
                 forvar43,
                 reg42,
                 reg40,
                 forvar39,
                 forvar38,
                 reg36,
                 reg35,
                 reg34,
                 reg32,
                 forvar31,
                 reg30,
                 forvar29,
                 forvar28,
                 (1'h0)};
  assign wire24 = wire21[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg25 <= ((((^(wire22 & wire20)) - wire21[(2'h3):(2'h3)]) ^~ (~&$unsigned($signed((8'ha0))))) & wire21[(1'h0):(1'h0)]);
    end
  assign wire26 = {$unsigned(wire22[(2'h2):(1'h1)])};
  always
    @(posedge clk) begin
      reg27 <= ($unsigned($signed(({wire22} ? {reg25, wire26} : wire23))) ?
          wire24 : wire24[(1'h1):(1'h0)]);
      for (forvar28 = (1'h0); (forvar28 < (2'h2)); forvar28 = (forvar28 + (1'h1)))
        begin
          for (forvar29 = (1'h0); (forvar29 < (3'h4)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 = wire21;
            end
          for (forvar31 = (1'h0); (forvar31 < (3'h4)); forvar31 = (forvar31 + (1'h1)))
            begin
              reg32 = "pmA5";
              reg33 <= $unsigned(reg27);
              reg34 = (&wire24[(3'h7):(3'h6)]);
              reg35 = $signed((&$signed(((forvar31 ? forvar29 : forvar29) ?
                  $signed(reg33) : (~^reg27)))));
            end
        end
      reg36 = $unsigned(wire20[(5'h10):(3'h4)]);
    end
  assign wire37 = reg27[(4'hd):(4'h8)];
  always
    @(posedge clk) begin
      for (forvar38 = (1'h0); (forvar38 < (3'h4)); forvar38 = (forvar38 + (1'h1)))
        begin
          for (forvar39 = (1'h0); (forvar39 < (3'h4)); forvar39 = (forvar39 + (1'h1)))
            begin
              reg40 = {wire24[(2'h3):(1'h0)], wire24[(1'h1):(1'h0)]};
              reg41 <= {($unsigned($unsigned($unsigned((8'ha1)))) ^ reg40)};
              reg42 = (wire20[(5'h14):(4'hf)] >> forvar38[(4'ha):(4'h9)]);
            end
        end
      for (forvar43 = (1'h0); (forvar43 < (3'h4)); forvar43 = (forvar43 + (1'h1)))
        begin
          for (forvar44 = (1'h0); (forvar44 < (2'h2)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 <= {wire26};
              reg46 = (forvar44 ^ wire24);
              reg47 <= ((~^{(+(~|(8'ha6))), wire20}) | reg45);
            end
          reg48 <= $signed((reg42 < reg42[(3'h5):(1'h1)]));
          reg49 <= (^~(8'hb0));
          for (forvar50 = (1'h0); (forvar50 < (1'h0)); forvar50 = (forvar50 + (1'h1)))
            begin
              reg51 <= $signed((((-wire22[(1'h1):(1'h1)]) ^ (~(reg48 >= forvar50))) ?
                  (|forvar44[(1'h0):(1'h0)]) : $unsigned(((reg47 != wire24) ?
                      (reg49 ? reg49 : wire37) : forvar39[(2'h3):(2'h2)]))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar52 = (1'h0); (forvar52 < (3'h4)); forvar52 = (forvar52 + (1'h1)))
        begin
          reg53 = (~|reg47[(2'h2):(1'h0)]);
          for (forvar54 = (1'h0); (forvar54 < (2'h3)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 <= $signed({$unsigned($signed($signed(reg49)))});
              reg56 = {wire26};
              reg57 <= $unsigned(($unsigned(reg33[(1'h1):(1'h1)]) ?
                  (reg55 + $signed((reg51 ?
                      reg49 : reg47))) : ($unsigned((reg47 ? reg33 : reg55)) ?
                      $unsigned((reg33 < wire20)) : ((reg47 ? reg56 : wire26) ?
                          (~^wire21) : (reg45 << reg49)))));
              reg58 = forvar52[(5'h12):(5'h11)];
              reg59 <= reg33;
            end
        end
    end
  assign wire60 = (({$unsigned((~^reg55)), reg57} ?
                          $signed({$unsigned(reg41),
                              {reg41,
                                  wire26}}) : $signed(reg57[(3'h7):(3'h4)])) ?
                      {{((reg33 || reg27) ?
                                  $signed(reg48) : reg27)}} : reg48[(3'h5):(3'h4)]);
  assign wire61 = $unsigned(reg57);
  always
    @(posedge clk) begin
      if ($unsigned($signed(reg47[(3'h5):(3'h5)])))
        begin
          reg62 <= ($signed(($signed((reg51 ? reg55 : reg45)) ?
                  $signed($signed(reg51)) : {$signed(reg25)})) ?
              $signed((~&reg45)) : (~^(~|{{reg47, wire20}})));
          reg63 = reg47[(1'h1):(1'h1)];
          reg64 <= (((^~(wire37 ~^ $signed(reg27))) ^ (wire60[(2'h3):(1'h1)] ?
                  ((reg62 > reg51) <= $unsigned(wire37)) : wire26[(3'h5):(2'h3)])) ?
              (|reg27[(4'he):(4'ha)]) : (8'hab));
        end
      else
        begin
          reg62 <= $signed(($signed(reg49[(3'h5):(1'h0)]) ?
              $unsigned((reg57[(3'h5):(2'h2)] | "K2po0P")) : $unsigned($signed(reg27))));
          for (forvar63 = (1'h0); (forvar63 < (1'h1)); forvar63 = (forvar63 + (1'h1)))
            begin
              reg64 <= (wire21[(3'h7):(3'h7)] ?
                  $unsigned((wire20[(3'h5):(2'h3)] << (reg48 << {(7'h40),
                      wire24}))) : wire37);
              reg65 <= wire60;
              reg66 = $unsigned(($signed((~&$signed(reg62))) >> reg59));
            end
          if (reg55[(1'h1):(1'h0)])
            begin
              reg67 <= (reg41 >> wire24[(3'h4):(3'h4)]);
              reg68 <= {wire24};
            end
          else
            begin
              reg67 <= $unsigned(wire37[(2'h2):(1'h0)]);
            end
        end
      reg69 = reg65[(4'h9):(1'h1)];
    end
  assign wire70 = ((~(~(wire21 ?
                      $unsigned((8'hba)) : reg47))) << ($unsigned(reg41[(4'h9):(2'h2)]) ?
                      reg41 : {{wire20}}));
  assign wire71 = $signed(((+$unsigned($unsigned(wire20))) ?
                      (wire61 ?
                          (reg67 ?
                              $unsigned((8'hb5)) : {reg25,
                                  wire22}) : {wire20[(5'h10):(3'h5)],
                              wire37[(3'h4):(2'h2)]}) : (wire26[(1'h1):(1'h0)] ?
                          (|reg59) : {(~reg25)})));
  always
    @(posedge clk) begin
      reg72 = (~|$unsigned(($signed(wire60[(4'ha):(2'h3)]) ?
          {wire61} : wire60[(2'h2):(1'h0)])));
      for (forvar73 = (1'h0); (forvar73 < (1'h0)); forvar73 = (forvar73 + (1'h1)))
        begin
          reg74 <= reg59;
          for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
            begin
              reg76 <= ((&($signed($signed(reg62)) ?
                      reg45 : {reg68[(3'h4):(2'h2)]})) ?
                  reg49 : {wire26});
              reg77 = $unsigned(reg55);
              reg78 = $unsigned(((&wire23[(1'h1):(1'h0)]) ?
                  {wire24[(3'h6):(2'h2)]} : $unsigned(wire37[(1'h1):(1'h1)])));
              reg79 <= reg45[(2'h3):(1'h0)];
            end
          reg80 <= {wire22, reg65};
          for (forvar81 = (1'h0); (forvar81 < (1'h1)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 <= reg62[(2'h2):(1'h0)];
            end
          for (forvar83 = (1'h0); (forvar83 < (1'h1)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 = reg80;
              reg85 <= forvar83[(3'h6):(3'h5)];
            end
        end
      if (wire71)
        begin
          for (forvar86 = (1'h0); (forvar86 < (1'h0)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 <= ({"cr7KS0W5Bngp",
                  $unsigned((forvar81 ?
                      $signed(reg27) : (8'h9f)))} * (-((wire61 ?
                  (wire37 != reg78) : reg33) || reg45[(2'h3):(2'h2)])));
              reg88 = wire26;
              reg89 <= {"8Puum", $unsigned(reg47)};
              reg90 = wire22;
              reg91 <= wire70[(2'h2):(1'h1)];
            end
          if ($unsigned($signed(($signed((wire23 ?
              reg62 : reg82)) << $unsigned((forvar83 && reg76))))))
            begin
              reg92 <= $unsigned((reg64 ? (8'hb4) : reg65[(4'hb):(2'h2)]));
              reg93 = $unsigned($signed((|((&reg55) ?
                  $signed(reg89) : $signed(reg59)))));
            end
          else
            begin
              reg92 <= forvar81[(3'h5):(2'h2)];
              reg94 <= wire21[(1'h1):(1'h0)];
              reg95 = (wire20 * (|$unsigned((wire23[(4'h8):(3'h4)] * (reg76 && wire61)))));
              reg96 = $signed((reg68 != (reg78 ?
                  reg74 : {reg51, $unsigned((8'hb2))})));
              reg97 <= (wire26 ?
                  (|$signed($signed((+forvar83)))) : (+(~&$signed(forvar75[(2'h2):(1'h0)]))));
            end
          reg98 = $signed(reg48);
        end
      else
        begin
          reg86 = $signed({reg76[(4'h8):(2'h2)]});
          reg87 <= $signed(((reg65 >> $signed((8'hb4))) ?
              ("g4" <= (^$signed(reg82))) : ((reg78[(2'h2):(1'h1)] * (+forvar81)) ?
                  (reg84 != (-wire22)) : (reg51 || (reg76 ? reg51 : reg48)))));
          reg88 = $unsigned(reg86[(3'h5):(3'h5)]);
        end
    end
endmodule
module top
#( parameter param810 = ((~^((~&(-(8'ha1))) ? (&(-(7'h44))) : {{(8'ha6), (7'h41)}, (^(8'ha2))})) ? ((((&(8'ha6)) ? ((8'h9f) ? (8'hbc) : (8'ha3)) : ((8'h9f) ? (8'ha4) : (8'ha0))) ? (((8'ha9) ? (8'hb1) : (8'h9e)) ? (!(8'ha7)) : ((8'ha2) ^ (8'hb0))) : (!((8'hb9) ? (7'h44) : (8'ha2)))) == (^(((7'h44) << (8'hae)) ^ ((7'h41) != (8'hba))))) : {((+((8'hb4) ? (8'hb0) : (8'hb3))) != (((8'hac) ? (8'hb8) : (8'ha7)) | ((8'ha0) >= (8'hbb)))), (+(((8'ha2) > (8'hb9)) << {(8'ha6)}))}) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h56d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire0;
  input wire signed [(5'h10):(1'h0)] wire1;
  input wire signed [(4'h8):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire3;
  input wire [(4'hd):(1'h0)] wire4;
  wire signed [(4'hb):(1'h0)] wire808;
  wire signed [(4'ha):(1'h0)] wire5;
  reg signed [(4'hb):(1'h0)] forvar6 = (1'h0);
  reg [(4'hb):(1'h0)] reg7 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar8 = (1'h0);
  reg signed [(4'he):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg10 = (1'h0);
  reg [(5'h10):(1'h0)] reg11 = (1'h0);
  reg [(4'hb):(1'h0)] reg12 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg [(4'hc):(1'h0)] reg14 = (1'h0);
  reg [(4'h9):(1'h0)] reg15 = (1'h0);
  reg [(4'h9):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg17 = (1'h0);
  reg [(4'he):(1'h0)] reg18 = (1'h0);
  reg [(3'h5):(1'h0)] reg19 = (1'h0);
  reg [(5'h13):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg82 = (1'h0);
  wire [(5'h11):(1'h0)] wire806;
  assign y = {wire808,
                 wire5,
                 forvar6,
                 reg7,
                 forvar8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg42,
                 reg82,
                 (1'h0)};
  assign wire5 = wire1;
  always
    @(posedge clk) begin
      for (forvar6 = (1'h0); (forvar6 < (2'h3)); forvar6 = (forvar6 + (1'h1)))
        begin
          reg7 = wire2;
          for (forvar8 = (1'h0); (forvar8 < (1'h0)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 = $signed({((^(wire0 >> wire0)) ?
                      $signed($unsigned((8'ha0))) : {reg7})});
            end
          reg10 = ($unsigned(wire1) <= wire0[(1'h0):(1'h0)]);
          reg11 = (~reg10);
        end
      if (wire1[(4'ha):(2'h2)])
        begin
          reg12 <= $unsigned(wire5[(3'h4):(1'h0)]);
          reg13 = $unsigned((+reg9));
          reg14 = $signed($signed((($unsigned(reg9) * $signed(wire1)) ?
              wire0[(2'h2):(1'h1)] : $signed($signed(wire2)))));
        end
      else
        begin
          if ($unsigned(({$unsigned((reg9 >>> wire1)), $signed($signed(reg9))} ?
              ((!reg12[(3'h7):(2'h2)]) ?
                  $signed("G38Y91HT") : reg12) : ($unsigned(reg7[(2'h2):(2'h2)]) ?
                  $signed($signed((8'ha6))) : {(reg9 * wire3),
                      forvar6[(3'h6):(2'h2)]}))))
            begin
              reg12 = $signed((reg9[(3'h6):(2'h2)] > (wire5 ? reg7 : reg12)));
              reg13 = $signed({{forvar6[(3'h4):(1'h0)]}});
            end
          reg15 <= wire2;
          reg16 = reg12[(4'ha):(3'h6)];
          if ((!{$unsigned($unsigned(wire4))}))
            begin
              reg17 <= $signed((($unsigned((wire1 ?
                      reg10 : wire1)) >>> (^{reg10})) ?
                  wire0 : wire4));
              reg18 <= reg12[(1'h0):(1'h0)];
              reg19 = (&reg11);
              reg42 <= $signed(((~&reg18[(4'hb):(3'h7)]) ?
                  (reg19 ?
                      (|(forvar6 ?
                          reg18 : (8'h9f))) : (wire1[(2'h3):(2'h3)] && $signed(reg12))) : (forvar6[(4'h9):(3'h4)] <= (+"CJTy"))));     
              reg82 = (!(8'hae));
            end
        end
    end
  module177 modinst807 (wire806, clk, reg9, reg11, wire4, reg42, reg82);
endmodule

module module177
#( parameter param804 = ((|({(~&(7'h40)), (^(7'h40))} ? {{(8'hb1), (8'hbe)}, {(8'hba), (8'ha8)}} : (8'hbb))) ? (|(~&(((7'h43) >= (8'hb8)) ? ((8'haa) | (8'h9e)) : ((8'hb4) & (8'hb7))))) : (~^(8'ha8)))
, parameter param805 = (&param804) )
(y, clk, wire178, wire179, wire180, wire181, wire182);
  output wire [(32'h307):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire178;
  input wire [(5'h10):(1'h0)] wire179;
  input wire [(4'hd):(1'h0)] wire180;
  input wire signed [(5'h13):(1'h0)] wire181;
  input wire signed [(4'hf):(1'h0)] wire182;
  wire [(2'h3):(1'h0)] wire183;
  reg signed [(4'he):(1'h0)] forvar184 = (1'h0);
  reg [(5'h14):(1'h0)] reg185 = (1'h0);
  reg signed [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(3'h4):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg [(5'h14):(1'h0)] reg189 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire190;
  wire signed [(5'h10):(1'h0)] wire191;
  wire [(5'h10):(1'h0)] wire192;
  wire [(4'h8):(1'h0)] wire347;
  wire signed [(4'hd):(1'h0)] wire451;
  assign y = {wire183,
                 forvar184,
                 reg185,
                 reg186,
                 reg187,
                 reg188,
                 reg189,
                 wire190,
                 wire191,
                 wire192,
                 wire347,
                 wire451,
                 (1'h0)};
  assign wire183 = ((^~(wire182[(2'h3):(2'h3)] == $signed("XtM2s3Eu"))) ?
                       wire182[(2'h3):(1'h1)] : $signed((8'hb8)));
  always
    @(posedge clk) begin
      for (forvar184 = (1'h0); (forvar184 < (3'h4)); forvar184 = (forvar184 + (1'h1)))
        begin
          reg185 = {(wire180 & (^((&wire183) ?
                  {forvar184, wire182} : forvar184[(4'h9):(2'h3)])))};
          reg186 = forvar184;
          reg187 <= wire179;
          reg188 = wire181[(1'h0):(1'h0)];
        end
      reg189 <= {wire178[(1'h0):(1'h0)], (|wire179[(2'h3):(1'h1)])};
    end
  assign wire191 = (~(!$signed(($unsigned(reg188) - reg187))));
  assign wire192 = $signed(wire179[(2'h3):(2'h2)]);
  module193 modinst348 (wire347, clk, reg189, wire192, wire179, reg188);
endmodule

module module193  (y, clk, wire197, wire196, wire195, wire194);
  output wire [(32'h6e4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire197;
  input wire signed [(5'h10):(1'h0)] wire196;
  input wire signed [(3'h6):(1'h0)] wire195;
  input wire [(4'hd):(1'h0)] wire194;
  reg signed [(5'h14):(1'h0)] reg204 = (1'h0);
  reg [(5'h15):(1'h0)] reg203 = (1'h0);
  reg [(5'h13):(1'h0)] reg202 = (1'h0);
  reg [(3'h7):(1'h0)] reg201 = (1'h0);
  reg [(4'hc):(1'h0)] forvar200 = (1'h0);
  reg [(5'h13):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar198 = (1'h0);
  assign y = {reg204,
                 reg203,
                 reg202,
                 reg201,
                 forvar200,
                 reg199,
                 forvar198,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar198 = (1'h0); (forvar198 < (1'h1)); forvar198 = (forvar198 + (1'h1)))
        begin
          reg199 = wire196[(3'h6):(3'h4)];
          for (forvar200 = (1'h0); (forvar200 < (2'h2)); forvar200 = (forvar200 + (1'h1)))
            begin
              reg201 = (&((^~$unsigned($signed(reg199))) ?
                  $unsigned(((^~forvar200) & (8'h9f))) : wire195));
              reg202 <= (~&$signed({($unsigned(forvar198) ?
                      $unsigned((7'h41)) : "5vXsSIrM"),
                  ("WCcbulRgPXMf3rRDI" ? "" : $unsigned(reg201))}));
              reg203 = (wire195[(1'h0):(1'h0)] == ((^~{$signed(reg199),
                      (wire196 ? reg199 : wire197)}) ?
                  (-$unsigned((^forvar200))) : (~^(reg202[(2'h3):(1'h0)] <<< $unsigned(wire197)))));
              reg204 <= $signed($unsigned($unsigned(wire196)));
            end
	end
    end
endmodule

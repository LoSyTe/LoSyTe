(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param774 = {(~(((|(8'hba)) ? {(8'hbf), (8'ha4)} : (|(7'h43))) ? (((7'h41) - (8'hbd)) ? ((7'h42) || (8'hac)) : (^~(8'had))) : (((8'ha2) ? (8'hbb) : (8'h9e)) ? ((8'hb3) > (8'h9f)) : ((8'hb6) <= (7'h40))))), ((~^((~(7'h40)) ? {(8'hbb)} : (~&(8'hb7)))) + (~&(((8'h9f) ? (8'h9d) : (8'ha4)) ? ((8'hac) >> (8'h9e)) : ((8'h9e) || (8'h9e)))))} )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h5d1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire0;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire signed [(4'hd):(1'h0)] wire3;
  wire [(4'h8):(1'h0)] wire773;
  wire signed [(5'h11):(1'h0)] wire772;
  reg [(5'h13):(1'h0)] reg771 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg768 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg767 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg766 = (1'h0);
  reg signed [(4'he):(1'h0)] reg765 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg764 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg763 = (1'h0);
  reg [(3'h4):(1'h0)] forvar762 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar761 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg760 = (1'h0);
  reg [(2'h3):(1'h0)] reg759 = (1'h0);
  reg [(4'ha):(1'h0)] reg758 = (1'h0);
  reg [(3'h4):(1'h0)] reg757 = (1'h0);
  reg [(4'hb):(1'h0)] forvar756 = (1'h0);
  reg [(5'h14):(1'h0)] forvar753 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg755 = (1'h0);
  reg [(2'h3):(1'h0)] reg754 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg753 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg752 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg751 = (1'h0);
  reg [(4'he):(1'h0)] reg750 = (1'h0);
  reg [(4'hd):(1'h0)] reg749 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg747 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg746 = (1'h0);
  reg [(4'h9):(1'h0)] reg745 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg744 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg743 = (1'h0);
  reg [(4'hf):(1'h0)] forvar742 = (1'h0);
  reg [(4'hd):(1'h0)] reg741 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire740;
  reg [(2'h3):(1'h0)] reg739 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg738 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg737 = (1'h0);
  reg [(4'he):(1'h0)] reg736 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar732 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg734 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg733 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg731 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg730 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg729 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg727 = (1'h0);
  reg [(5'h13):(1'h0)] reg726 = (1'h0);
  reg [(4'h8):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg724 = (1'h0);
  reg [(4'hf):(1'h0)] forvar720 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg723 = (1'h0);
  reg signed [(4'he):(1'h0)] reg722 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg721 = (1'h0);
  reg [(4'h8):(1'h0)] reg720 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire719;
  reg [(4'he):(1'h0)] reg718 = (1'h0);
  reg [(5'h13):(1'h0)] reg717 = (1'h0);
  reg [(5'h13):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg714 = (1'h0);
  reg [(4'ha):(1'h0)] reg713 = (1'h0);
  reg [(3'h4):(1'h0)] reg712 = (1'h0);
  reg [(4'he):(1'h0)] reg711 = (1'h0);
  reg [(4'hd):(1'h0)] reg710 = (1'h0);
  reg [(4'he):(1'h0)] reg709 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg708 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar707 = (1'h0);
  reg [(5'h13):(1'h0)] reg706 = (1'h0);
  reg [(5'h13):(1'h0)] reg705 = (1'h0);
  reg [(2'h3):(1'h0)] reg704 = (1'h0);
  reg [(3'h7):(1'h0)] reg703 = (1'h0);
  reg [(5'h10):(1'h0)] reg702 = (1'h0);
  reg [(3'h5):(1'h0)] forvar701 = (1'h0);
  reg [(2'h3):(1'h0)] reg700 = (1'h0);
  reg [(4'he):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg697 = (1'h0);
  reg [(2'h3):(1'h0)] forvar696 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg695 = (1'h0);
  reg [(4'h9):(1'h0)] reg694 = (1'h0);
  reg [(4'hf):(1'h0)] reg693 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar688 = (1'h0);
  reg [(5'h15):(1'h0)] reg692 = (1'h0);
  reg [(4'hb):(1'h0)] reg691 = (1'h0);
  reg [(4'ha):(1'h0)] forvar690 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg688 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg687 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg686 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg685 = (1'h0);
  reg [(3'h7):(1'h0)] reg684 = (1'h0);
  reg [(5'h14):(1'h0)] reg683 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar682 = (1'h0);
  reg [(3'h7):(1'h0)] forvar681 = (1'h0);
  reg [(2'h3):(1'h0)] reg680 = (1'h0);
  reg [(3'h7):(1'h0)] reg679 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire678;
  wire signed [(4'h9):(1'h0)] wire676;
  wire [(2'h2):(1'h0)] wire675;
  wire [(4'hc):(1'h0)] wire674;
  reg [(5'h12):(1'h0)] reg4 = (1'h0);
  reg [(5'h15):(1'h0)] forvar5 = (1'h0);
  reg [(4'hb):(1'h0)] reg6 = (1'h0);
  reg [(4'h8):(1'h0)] reg7 = (1'h0);
  reg [(4'h8):(1'h0)] reg8 = (1'h0);
  reg [(5'h12):(1'h0)] forvar9 = (1'h0);
  reg [(5'h11):(1'h0)] reg10 = (1'h0);
  reg [(3'h6):(1'h0)] reg11 = (1'h0);
  reg signed [(4'he):(1'h0)] reg12 = (1'h0);
  reg [(5'h12):(1'h0)] reg13 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg14 = (1'h0);
  reg [(5'h10):(1'h0)] reg9 = (1'h0);
  reg [(5'h12):(1'h0)] reg15 = (1'h0);
  reg [(4'ha):(1'h0)] forvar16 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg17 = (1'h0);
  reg [(3'h5):(1'h0)] forvar18 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg19 = (1'h0);
  reg [(5'h15):(1'h0)] forvar20 = (1'h0);
  reg [(4'hb):(1'h0)] reg21 = (1'h0);
  wire [(3'h4):(1'h0)] wire669;
  wire [(5'h11):(1'h0)] wire671;
  wire [(5'h10):(1'h0)] wire672;
  assign y = {wire773,
                 wire772,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 reg765,
                 reg764,
                 reg763,
                 forvar762,
                 forvar761,
                 reg760,
                 reg759,
                 reg758,
                 reg757,
                 forvar756,
                 forvar753,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 forvar748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 forvar742,
                 reg741,
                 wire740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 forvar732,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 forvar720,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 wire719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 forvar707,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 forvar701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 forvar696,
                 reg695,
                 reg694,
                 reg693,
                 reg690,
                 forvar688,
                 reg692,
                 reg691,
                 forvar690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 forvar682,
                 forvar681,
                 reg680,
                 reg679,
                 wire678,
                 wire676,
                 wire675,
                 wire674,
                 reg4,
                 forvar5,
                 reg6,
                 reg7,
                 reg8,
                 forvar9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg9,
                 reg15,
                 forvar16,
                 reg17,
                 forvar18,
                 reg19,
                 forvar20,
                 reg21,
                 wire669,
                 wire671,
                 wire672,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 = wire1[(3'h4):(3'h4)];
      if ({((^~(^$signed(reg4))) * wire2)})
        begin
          for (forvar5 = (1'h0); (forvar5 < (2'h2)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg6 <= (~|((~|{$signed(wire2), wire2}) && forvar5));
              reg7 = $unsigned(wire2);
            end
          reg8 <= (8'hb2);
          for (forvar9 = (1'h0); (forvar9 < (1'h0)); forvar9 = (forvar9 + (1'h1)))
            begin
              reg10 <= wire1;
              reg11 <= wire2[(4'hc):(4'h9)];
              reg12 <= ({$unsigned($signed((&reg11)))} ?
                  wire0[(4'hc):(3'h4)] : {$unsigned($signed(forvar5)),
                      (~^wire3[(1'h0):(1'h0)])});
              reg13 <= $signed($signed(wire2));
            end
          reg14 <= (((!((-forvar5) ?
                  wire0 : $signed(wire3))) | $unsigned({$unsigned(reg12)})) ?
              $signed($signed(wire2)) : $unsigned((-wire0[(4'ha):(3'h7)])));
        end
      else
        begin
          for (forvar5 = (1'h0); (forvar5 < (1'h0)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg6 = (&({$unsigned(reg13), (((8'haf) >>> wire1) - {reg11})} ?
                  $unsigned(wire2[(4'ha):(3'h5)]) : $signed($unsigned((reg12 ?
                      (8'hb8) : reg7)))));
              reg7 <= ($signed(reg11[(1'h0):(1'h0)]) * reg7);
              reg8 = $unsigned((~reg12));
              reg9 <= $unsigned(wire2);
              reg10 = forvar5[(5'h14):(5'h13)];
            end
          if (((((|$unsigned((8'hb4))) <<< ((reg6 ?
                  (8'hb8) : (8'had)) << $unsigned(wire3))) ?
              $signed($unsigned($signed(reg6))) : $unsigned($signed($unsigned(reg9)))) <<< {forvar9,
              (~^reg11)}))
            begin
              reg11 = $signed(((7'h44) ?
                  wire2[(4'hc):(1'h0)] : $signed($unsigned(((8'ha2) ?
                      reg8 : (8'had))))));
              reg12 <= (reg8 ? (^wire3) : wire1);
            end
          else
            begin
              reg11 = ((forvar5 > forvar5[(4'h9):(2'h3)]) ?
                  reg11 : (~reg11[(1'h1):(1'h1)]));
              reg12 <= reg13[(4'hb):(3'h5)];
              reg13 <= $signed($signed($signed({(reg8 ? forvar9 : wire1)})));
              reg14 <= (!wire1);
            end
          reg15 = ((wire2 ^ {reg12[(2'h2):(1'h0)]}) && $signed($signed({(wire0 ?
                  forvar5 : reg12),
              reg11})));
        end
      for (forvar16 = (1'h0); (forvar16 < (1'h0)); forvar16 = (forvar16 + (1'h1)))
        begin
          reg17 <= $unsigned(($signed($unsigned($unsigned(reg8))) || forvar5[(4'hb):(3'h4)]));
          for (forvar18 = (1'h0); (forvar18 < (3'h4)); forvar18 = (forvar18 + (1'h1)))
            begin
              reg19 <= $unsigned(reg11);
            end
        end
      for (forvar20 = (1'h0); (forvar20 < (1'h0)); forvar20 = (forvar20 + (1'h1)))
        begin
          reg21 <= $unsigned(($unsigned($unsigned($signed(reg9))) ?
              $unsigned((~&reg4)) : forvar16));
        end
    end
  module22 modinst670 (.wire23(forvar20), .wire25(wire2), .y(wire669), .wire26(reg4), .wire24(reg15), .clk(clk));
  assign wire671 = {((~^{(reg10 ~^ reg17), {forvar16}}) ?
                           reg6[(3'h4):(1'h1)] : (|(~&((8'hbd) ^~ reg8))))};
  module412 modinst673 (wire672, clk, reg12, forvar9, wire671, reg19, reg15);
  assign wire674 = (|"4uqDSd");
  assign wire675 = wire672;
  module29 modinst677 (.wire32(wire674), .clk(clk), .wire30(wire672), .wire33(wire2), .y(wire676), .wire31(reg13));
  assign wire678 = reg12[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg679 <= $unsigned(reg6[(4'h8):(1'h0)]);
      reg680 = reg679[(2'h3):(2'h2)];
      for (forvar681 = (1'h0); (forvar681 < (3'h4)); forvar681 = (forvar681 + (1'h1)))
        begin
          for (forvar682 = (1'h0); (forvar682 < (2'h3)); forvar682 = (forvar682 + (1'h1)))
            begin
              reg683 <= $signed(wire672[(4'hc):(4'h8)]);
              reg684 = forvar18;
              reg685 = ({{(^~((8'hb1) && reg15))}} ?
                  (~^{reg14[(4'h8):(3'h7)]}) : (!((reg6[(4'h8):(3'h7)] ?
                      reg8 : {(8'hae)}) >= wire672[(4'hc):(3'h5)])));
              reg686 = ((~|wire678) ?
                  (~&$signed({wire672,
                      (~&reg8)})) : ($signed($unsigned($signed((8'hb4)))) & $unsigned($unsigned((wire675 ?
                      reg685 : wire1)))));
            end
        end
      reg687 = (~&(reg21 ?
          reg685 : (($signed(reg4) && ((8'ha9) ? (7'h43) : forvar18)) ?
              wire0[(3'h7):(3'h4)] : $unsigned(reg6[(3'h5):(2'h3)]))));
      if ((($unsigned((~&{wire675, wire0})) - ($signed({reg687,
              wire3}) >>> wire676[(4'h8):(1'h1)])) ?
          {$unsigned((!(wire674 >>> (8'had)))),
              "Fmz293DYEkJ"} : {((|(reg4 | reg680)) ?
                  (wire1 & (~|(8'hbc))) : $signed($unsigned(wire671)))}))
        begin
          reg688 <= wire2;
          if ($unsigned((~reg684)))
            begin
              reg689 = ({forvar681} ?
                  ("BHhomT" || reg680[(1'h0):(1'h0)]) : $signed($unsigned(reg684)));
            end
          else
            begin
              reg689 <= $signed(($unsigned(reg17) ?
                  $signed($signed(((8'hba) ^~ (8'ha8)))) : ($unsigned(forvar16) ?
                      {(reg11 <<< forvar5),
                          (forvar9 ^~ forvar5)} : (reg7[(3'h6):(2'h2)] ?
                          (forvar9 == reg9) : (8'hb7)))));
            end
          for (forvar690 = (1'h0); (forvar690 < (1'h1)); forvar690 = (forvar690 + (1'h1)))
            begin
              reg691 <= $signed(forvar20);
            end
          reg692 <= (-"acBSqQLHG7E7GhRoYOKo");
        end
      else
        begin
          for (forvar688 = (1'h0); (forvar688 < (1'h1)); forvar688 = (forvar688 + (1'h1)))
            begin
              reg689 <= wire2[(3'h4):(2'h2)];
              reg690 <= (^(^"eln0ml3QCg2c5v5"));
            end
          if (($signed({$unsigned(reg680),
              $unsigned(wire678)}) <<< reg13[(4'hf):(4'ha)]))
            begin
              reg691 = wire2[(4'hb):(3'h5)];
            end
          else
            begin
              reg691 <= $unsigned({{(reg10 ?
                          (forvar682 < reg683) : $signed((8'ha5))),
                      $unsigned((^~forvar5))}});
              reg692 <= $signed(((($signed(reg679) ?
                          {reg17, reg7} : reg13[(1'h0):(1'h0)]) ?
                      $unsigned((^reg6)) : forvar688) ?
                  $unsigned(reg4[(4'h8):(3'h6)]) : reg9[(4'hf):(1'h0)]));
              reg693 <= $unsigned($unsigned(reg692));
              reg694 = wire0[(4'hd):(3'h4)];
              reg695 <= reg685[(3'h4):(2'h3)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar696 = (1'h0); (forvar696 < (2'h2)); forvar696 = (forvar696 + (1'h1)))
        begin
          if (($unsigned(({$signed(reg8)} ?
                  reg693[(4'he):(4'hc)] : $unsigned($unsigned((8'haf))))) ?
              (~^forvar20[(3'h5):(3'h5)]) : (!{(+(^(8'ha3)))})))
            begin
              reg697 <= (reg4 ^ ((^$signed((~^reg7))) ~^ ({$unsigned(reg690)} + $signed((8'ha8)))));
            end
          else
            begin
              reg697 <= {{(8'hbb)}, reg684[(3'h7):(2'h2)]};
              reg698 = (~|reg21);
              reg699 = ($signed(wire676[(2'h3):(2'h3)]) ?
                  $unsigned((^~$unsigned(reg690[(3'h6):(2'h3)]))) : $signed((reg15 >= ($unsigned(forvar688) | $signed(wire0)))));
              reg700 = $unsigned({(^{(~&wire669),
                      (reg698 ? reg685 : reg680)})});
            end
          for (forvar701 = (1'h0); (forvar701 < (3'h4)); forvar701 = (forvar701 + (1'h1)))
            begin
              reg702 <= (((reg691[(3'h5):(3'h4)] | (&{forvar696,
                      reg695})) >= (($signed(forvar18) ?
                          (wire1 ? (8'hb9) : forvar701) : reg688) ?
                      reg689[(4'hf):(1'h1)] : $unsigned(forvar9))) ?
                  $signed($signed(((|forvar5) <= $unsigned(wire3)))) : ((+reg6[(4'ha):(3'h7)]) ?
                      $signed(reg8) : (~&(~^(reg700 ? (8'hbf) : forvar701)))));
              reg703 <= (($signed(($signed((8'ha6)) * (reg4 <<< reg7))) ^ (~^reg692)) ?
                  wire3 : reg15);
              reg704 = ({reg694[(2'h2):(1'h0)],
                  $unsigned(wire675[(1'h1):(1'h1)])} & reg12[(3'h7):(3'h4)]);
              reg705 <= (reg13[(1'h1):(1'h0)] < ((({reg679} || (8'hbc)) ^~ (~&$signed(reg684))) ?
                  $signed(($unsigned(reg6) ?
                      $unsigned(forvar690) : reg14[(3'h4):(1'h0)])) : $unsigned((~&$signed(reg19)))));
              reg706 <= ($unsigned($unsigned($signed((^(8'ha5))))) * wire2);
            end
        end
      for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
        begin
          if ($unsigned((^(reg695 + (~^(forvar688 ^ reg698))))))
            begin
              reg708 <= $signed(wire674[(3'h4):(2'h3)]);
              reg709 = forvar9;
              reg710 <= forvar9[(3'h7):(1'h0)];
              reg711 = reg691;
            end
          else
            begin
              reg708 <= reg711;
            end
          if (((reg19 | (^(+(+forvar701)))) ?
              ($unsigned(({wire2, wire672} ?
                  (wire678 ?
                      forvar18 : reg691) : ((8'hae) >= reg698))) <<< (!$signed((forvar701 ?
                  reg711 : reg698)))) : ($signed(($signed((7'h44)) < $signed(reg705))) > reg690[(4'hb):(4'ha)])))
            begin
              reg712 <= (reg710[(3'h6):(1'h1)] != reg10[(4'ha):(2'h3)]);
              reg713 = "2FRFckLphAqYJm";
              reg714 <= ($unsigned(reg699) ?
                  $unsigned((+{$signed(reg9)})) : $signed(($unsigned($signed((8'haf))) ^~ {(~&forvar696),
                      ""})));
              reg715 <= ($signed(($signed((forvar696 && reg688)) - $signed({(8'h9c),
                      (8'ha0)}))) ?
                  $signed(forvar5) : {(~^(reg702[(4'he):(3'h7)] <<< (wire3 ?
                          reg704 : reg692))),
                      $signed(((8'hb3) ^~ reg708[(2'h2):(2'h2)]))});
              reg716 <= reg683[(4'hd):(2'h3)];
            end
          else
            begin
              reg712 <= (8'hb9);
              reg713 = ((wire671[(2'h3):(2'h2)] >>> ({(reg697 + reg716)} ?
                  reg680[(1'h0):(1'h0)] : ((reg689 << reg19) ?
                      (^~reg691) : $unsigned(reg691)))) ^~ $signed($unsigned(($unsigned(reg690) || reg695))));
              reg714 <= reg14;
            end
          reg717 = (reg714[(3'h5):(2'h2)] ?
              reg688[(4'hf):(3'h6)] : (reg4[(4'hf):(1'h1)] <<< ({(8'hb9),
                      (reg689 * reg692)} ?
                  ((reg691 ? forvar18 : wire674) ?
                      $signed(reg703) : (reg17 ?
                          reg686 : reg699)) : (-(wire675 ? reg13 : reg7)))));
          reg718 = reg716;
        end
    end
  assign wire719 = reg17[(4'hd):(2'h3)];
  always
    @(posedge clk) begin
      if ($signed($signed($unsigned($signed(reg685[(3'h6):(3'h4)])))))
        begin
          if ($unsigned(((forvar690[(1'h0):(1'h0)] ?
                  {(wire0 ? (7'h42) : reg688)} : $unsigned("96t3l")) ?
              reg7 : $signed("QD"))))
            begin
              reg720 <= ((reg686 ?
                      $unsigned("Y") : ($unsigned(reg709) ?
                          $unsigned(reg6[(3'h5):(2'h2)]) : ((~|reg712) ?
                              $signed(reg708) : (wire2 == reg12)))) ?
                  reg15[(5'h11):(1'h0)] : $unsigned((($signed(reg7) >= reg684[(3'h4):(3'h4)]) ?
                      ($unsigned(forvar690) * {forvar688}) : reg11)));
              reg721 <= (|$unsigned("YufbJOknkX484pqIG1v"));
            end
          else
            begin
              reg720 <= (8'h9d);
              reg721 <= wire675;
              reg722 <= $unsigned((&{(!wire672[(4'ha):(1'h1)]),
                  $signed((reg718 == wire3))}));
              reg723 <= reg708[(2'h3):(1'h1)];
            end
        end
      else
        begin
          for (forvar720 = (1'h0); (forvar720 < (1'h0)); forvar720 = (forvar720 + (1'h1)))
            begin
              reg721 = $unsigned((&$unsigned($unsigned((reg686 == reg691)))));
              reg722 <= ({reg709} >> $unsigned(($unsigned(reg694) || (((8'had) >>> wire2) + {reg683}))));
              reg723 <= reg7;
              reg724 <= ((~^(-((&wire3) ?
                  ((7'h44) ? forvar9 : reg721) : (reg694 ?
                      reg708 : (8'hb3))))) >= reg706);
              reg725 <= ($unsigned(reg680) ?
                  $signed($unsigned($unsigned($unsigned(reg724)))) : {$signed(forvar688[(4'hb):(2'h2)]),
                      ($signed(forvar701[(1'h0):(1'h0)]) ?
                          (^$signed(forvar696)) : forvar9[(4'he):(4'ha)])});
            end
          if ($signed($unsigned(wire678)))
            begin
              reg726 <= {{$signed($signed(reg690[(2'h2):(2'h2)]))},
                  $signed((+(wire672[(1'h1):(1'h0)] ?
                      "ythKgWFRYpDhIMF616" : reg723)))};
              reg727 <= $signed((forvar696 + ({$unsigned(reg703), {reg703}} ?
                  reg4[(3'h5):(2'h3)] : ((8'h9e) == (reg687 ?
                      reg12 : reg705)))));
            end
          else
            begin
              reg726 <= $signed($unsigned($signed(reg15[(4'ha):(3'h4)])));
              reg727 <= {(-{forvar707[(1'h0):(1'h0)]}), reg723};
              reg728 = $signed($unsigned(({((8'hb1) ~^ reg684)} ?
                  $signed("e1urVI") : wire672[(4'ha):(3'h5)])));
              reg729 <= (~$unsigned(($unsigned({reg722,
                  reg13}) ^ (reg693[(4'h8):(2'h2)] == (^~reg714)))));
              reg730 = wire2[(4'he):(4'h9)];
            end
        end
      if ((&wire674[(4'ha):(2'h2)]))
        begin
          if ($unsigned((-($signed((wire0 ?
              reg711 : reg680)) && (reg14[(3'h5):(3'h4)] ?
              reg712[(2'h3):(1'h1)] : (|wire3))))))
            begin
              reg731 <= {(-(~|({wire672} ?
                      forvar707[(3'h4):(1'h1)] : (reg14 >= (8'hba))))),
                  ((8'ha5) ?
                      (!(+$unsigned((8'ha8)))) : $unsigned(reg690[(1'h0):(1'h0)]))};
            end
          else
            begin
              reg731 <= forvar707;
              reg732 <= (~(($unsigned(reg716) ? reg19 : (^$unsigned(wire676))) ?
                  $signed(($unsigned(forvar688) ^ (7'h44))) : forvar707));
              reg733 = reg699;
              reg734 <= {$signed((($unsigned(reg704) ?
                          (reg706 ? reg10 : wire674) : $signed(wire669)) ?
                      ("ZLFvvsMvcXS" + forvar16) : (~|{reg722, reg723}))),
                  $signed(((+$unsigned(reg7)) >>> (-wire676)))};
            end
        end
      else
        begin
          reg731 = (wire1 ?
              $signed($signed((-reg717))) : (reg688 ?
                  reg14[(2'h2):(1'h1)] : $signed({reg716,
                      reg9[(3'h5):(3'h4)]})));
          for (forvar732 = (1'h0); (forvar732 < (2'h3)); forvar732 = (forvar732 + (1'h1)))
            begin
              reg733 <= "WW";
              reg734 = (($unsigned($unsigned(((8'ha9) ?
                  reg684 : wire672))) ^ wire672) | (!reg679[(1'h1):(1'h0)]));
              reg735 <= $unsigned($unsigned($unsigned($unsigned($signed((7'h44))))));
              reg736 = reg689[(5'h11):(4'hb)];
              reg737 = (reg711 ?
                  reg706 : $unsigned($signed(forvar690[(4'h9):(3'h6)])));
            end
        end
      reg738 <= $signed(({((forvar20 > reg686) ?
              (reg703 ?
                  reg702 : (8'ha0)) : $unsigned(wire674))} >>> reg729[(3'h7):(2'h2)]));
      reg739 <= (^~{reg736[(1'h1):(1'h0)]});
    end
  assign wire740 = (({(8'hb0),
                       ((forvar5 <= reg724) > $unsigned((8'ha3)))} <= forvar732[(4'h8):(3'h6)]) - $signed($unsigned(forvar688[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      if ((reg698 ? reg734 : $unsigned(forvar5[(4'hc):(4'h9)])))
        begin
          reg741 <= {(|(!reg685[(2'h2):(2'h2)]))};
          for (forvar742 = (1'h0); (forvar742 < (2'h2)); forvar742 = (forvar742 + (1'h1)))
            begin
              reg743 <= (^~({("rfB6" >>> (wire678 ? reg741 : reg697)),
                  $signed({reg687})} >> reg728));
              reg744 <= (reg6 != (reg737 ?
                  (&((wire0 >> reg704) + $signed(reg17))) : $signed($unsigned($unsigned(forvar720)))));
              reg745 <= $signed({(reg725[(3'h5):(1'h1)] ?
                      $signed(reg706) : (reg728[(3'h7):(1'h0)] ?
                          $unsigned(forvar18) : $signed(wire1)))});
              reg746 = reg6[(4'h9):(2'h3)];
              reg747 = reg13;
            end
          for (forvar748 = (1'h0); (forvar748 < (2'h3)); forvar748 = (forvar748 + (1'h1)))
            begin
              reg749 <= $unsigned($unsigned(($unsigned(reg747) > $signed((reg686 ?
                  reg697 : reg692)))));
              reg750 = (reg15[(1'h0):(1'h0)] & ((reg695[(2'h3):(1'h1)] ?
                  $signed({reg726,
                      wire2}) : $signed($signed(reg736))) <<< reg697[(2'h2):(1'h1)]));
              reg751 <= $unsigned({reg10});
              reg752 <= (~&{{(-forvar682[(3'h7):(3'h4)]),
                      ((reg695 || wire740) ? reg712 : forvar742)},
                  (wire0 < {(reg728 && (8'hba))})});
            end
        end
      else
        begin
          reg741 <= reg747[(2'h3):(1'h1)];
          for (forvar742 = (1'h0); (forvar742 < (3'h4)); forvar742 = (forvar742 + (1'h1)))
            begin
              reg743 <= reg21;
              reg744 <= (^~(!(&((&reg739) ^ reg698))));
              reg745 = reg732[(4'hc):(3'h5)];
              reg746 <= ((8'haa) ? (|reg710) : (~|reg697[(4'h8):(3'h6)]));
              reg747 <= (reg717[(5'h12):(4'hd)] & $signed((($signed(reg688) ?
                      (reg691 >= reg13) : (reg4 & (8'hac))) ?
                  ((reg724 || wire671) ?
                      (forvar742 ?
                          forvar20 : wire1) : $unsigned(reg699)) : {((8'hb3) ?
                          reg735 : (8'hae)),
                      ((8'h9e) == reg13)})));
            end
        end
      if ((-(+reg712[(1'h1):(1'h0)])))
        begin
          if (($signed(reg733[(3'h4):(3'h4)]) ~^ ($unsigned((reg727[(4'ha):(2'h2)] >= reg727)) ?
              reg13 : $unsigned($signed(reg700)))))
            begin
              reg753 = (({(&(8'ha5))} >> reg11[(3'h4):(1'h1)]) == "oNilhscJrmZgD57hNY2t");
              reg754 <= (8'ha2);
              reg755 <= $signed({(~&((wire2 ?
                      forvar682 : (8'ha8)) != reg726))});
            end
          else
            begin
              reg753 <= $signed($signed(reg685));
              reg754 <= wire671;
            end
        end
      else
        begin
          for (forvar753 = (1'h0); (forvar753 < (1'h1)); forvar753 = (forvar753 + (1'h1)))
            begin
              reg754 <= reg749[(4'hd):(3'h6)];
              reg755 <= $signed((reg705[(4'hd):(1'h0)] + {reg728,
                  {(~|reg746)}}));
            end
          for (forvar756 = (1'h0); (forvar756 < (2'h2)); forvar756 = (forvar756 + (1'h1)))
            begin
              reg757 <= "tb3xyTSMk7Bd";
              reg758 = "2liUnZGLVT44";
            end
        end
      reg759 = $unsigned(wire719[(2'h3):(1'h1)]);
      reg760 <= (reg749[(3'h4):(2'h2)] || reg732);
      for (forvar761 = (1'h0); (forvar761 < (1'h0)); forvar761 = (forvar761 + (1'h1)))
        begin
          for (forvar762 = (1'h0); (forvar762 < (3'h4)); forvar762 = (forvar762 + (1'h1)))
            begin
              reg763 <= reg743;
              reg764 = forvar682[(2'h3):(1'h1)];
            end
          reg765 <= reg6;
          reg766 <= "Dpaz4NrYnSRTMvIdh";
          if ($signed(reg735[(4'hc):(3'h6)]))
            begin
              reg767 <= ((7'h41) ?
                  $unsigned(reg11[(2'h3):(2'h3)]) : ($unsigned($signed((reg688 ?
                          wire3 : wire3))) ?
                      reg741[(3'h5):(2'h3)] : reg753[(3'h5):(2'h3)]));
              reg768 <= (^reg706);
              reg769 <= (&reg758[(3'h7):(3'h5)]);
            end
          else
            begin
              reg767 = reg686[(1'h0):(1'h0)];
              reg768 <= $signed($signed(reg693));
              reg769 <= ((forvar707 ~^ (reg750[(2'h2):(1'h1)] & (^~((7'h41) ?
                      reg752 : reg745)))) ?
                  forvar696[(1'h1):(1'h1)] : reg715);
              reg770 = ((reg741[(2'h2):(2'h2)] ?
                      $signed(((forvar9 ?
                          reg726 : wire740) - (!reg721))) : (($unsigned(reg19) ?
                          (-(7'h43)) : reg17[(4'hf):(1'h0)]) ^ $signed(((8'hb7) ?
                          reg700 : reg19)))) ?
                  $unsigned(reg692[(3'h5):(3'h5)]) : (8'hba));
              reg771 <= ($signed({(reg755[(3'h4):(3'h4)] + "VwKLJymMZOFgFDbG1KWK"),
                      (&wire671[(3'h4):(1'h1)])}) ?
                  (~^($signed(reg693[(4'hb):(3'h5)]) << (~^wire719[(2'h3):(1'h0)]))) : $signed($signed(reg736[(3'h6):(3'h5)])));
            end
        end
    end
  assign wire772 = (reg726[(3'h7):(2'h2)] ?
                       ((~$signed(reg770[(3'h6):(1'h1)])) ?
                           (reg725 ?
                               ((~(8'hb4)) ?
                                   $signed(reg12) : reg709) : $signed((!reg731))) : (~$unsigned($signed((8'ha3))))) : $unsigned(reg765[(1'h0):(1'h0)]));
  assign wire773 = reg757;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module22
#( parameter param668 = (((+(^~((8'ha8) ? (7'h42) : (8'hba)))) + (({(8'haa), (8'had)} + ((8'hb6) ? (7'h40) : (7'h40))) ? ({(8'hb6)} >> (|(8'hbe))) : ((~|(8'hb7)) <<< {(8'hb0), (8'hae)}))) | ({{((8'haf) >> (8'hb9))}} ? ((((8'h9c) ? (8'haa) : (8'hae)) ? ((8'ha1) <= (8'ha4)) : ((8'h9d) && (8'ha8))) > ((^~(8'hab)) < (~^(8'hb2)))) : (({(8'hb4)} ? ((8'ha7) ? (8'ha1) : (8'ha6)) : {(8'haf)}) ? (((8'hbd) ? (8'haf) : (8'hb4)) ? ((8'hae) ? (7'h43) : (8'hb1)) : (~^(8'hb4))) : (~^((8'had) <= (8'ha1)))))) )
(y, clk, wire26, wire25, wire24, wire23);
  output wire [(32'h643):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire26;
  input wire signed [(5'h14):(1'h0)] wire25;
  input wire signed [(2'h2):(1'h0)] wire24;
  input wire signed [(5'h15):(1'h0)] wire23;
  reg signed [(4'hf):(1'h0)] reg667 = (1'h0);
  reg [(4'ha):(1'h0)] forvar659 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg658 = (1'h0);
  reg [(2'h3):(1'h0)] reg666 = (1'h0);
  reg signed [(4'he):(1'h0)] reg665 = (1'h0);
  reg [(3'h4):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg663 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg662 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg661 = (1'h0);
  reg [(5'h14):(1'h0)] reg660 = (1'h0);
  reg [(5'h15):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar658 = (1'h0);
  reg [(4'ha):(1'h0)] reg657 = (1'h0);
  reg [(5'h10):(1'h0)] reg656 = (1'h0);
  reg [(4'h9):(1'h0)] reg655 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg654 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg653 = (1'h0);
  reg [(5'h12):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar651 = (1'h0);
  reg [(4'hb):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg648 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar647 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg646 = (1'h0);
  reg [(4'hc):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar642 = (1'h0);
  reg [(4'hc):(1'h0)] reg641 = (1'h0);
  reg [(5'h10):(1'h0)] forvar640 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire639;
  reg signed [(5'h12):(1'h0)] reg638 = (1'h0);
  reg [(3'h4):(1'h0)] reg637 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar636 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg635 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg633 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg631 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar630 = (1'h0);
  reg [(4'he):(1'h0)] reg629 = (1'h0);
  reg [(4'ha):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg627 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar626 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar624 = (1'h0);
  reg [(4'hb):(1'h0)] reg623 = (1'h0);
  reg [(4'h9):(1'h0)] reg622 = (1'h0);
  reg [(3'h6):(1'h0)] reg621 = (1'h0);
  reg [(2'h2):(1'h0)] reg620 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg619 = (1'h0);
  reg [(3'h4):(1'h0)] forvar618 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg617 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg615 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg614 = (1'h0);
  reg [(5'h11):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar612 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg611 = (1'h0);
  reg [(2'h3):(1'h0)] reg610 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg609 = (1'h0);
  reg [(3'h7):(1'h0)] reg608 = (1'h0);
  reg [(4'hd):(1'h0)] reg607 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg606 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar605 = (1'h0);
  reg [(4'ha):(1'h0)] reg604 = (1'h0);
  reg [(4'hd):(1'h0)] reg603 = (1'h0);
  reg [(4'he):(1'h0)] reg602 = (1'h0);
  reg [(2'h3):(1'h0)] reg601 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg600 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar599 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar598 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire597;
  reg [(4'h9):(1'h0)] reg596 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg595 = (1'h0);
  reg [(5'h13):(1'h0)] reg594 = (1'h0);
  reg [(4'hf):(1'h0)] forvar593 = (1'h0);
  reg [(4'he):(1'h0)] reg592 = (1'h0);
  reg [(5'h15):(1'h0)] reg591 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg590 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg589 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg588 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar587 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar585 = (1'h0);
  reg [(3'h5):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg583 = (1'h0);
  reg [(3'h5):(1'h0)] reg582 = (1'h0);
  reg [(4'ha):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg580 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar579 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg578 = (1'h0);
  reg [(3'h4):(1'h0)] reg577 = (1'h0);
  reg [(5'h15):(1'h0)] reg576 = (1'h0);
  reg [(4'hd):(1'h0)] forvar575 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg573 = (1'h0);
  wire [(4'he):(1'h0)] wire572;
  wire [(3'h6):(1'h0)] wire567;
  wire signed [(5'h13):(1'h0)] wire566;
  wire signed [(5'h15):(1'h0)] wire565;
  wire signed [(3'h6):(1'h0)] wire561;
  wire signed [(4'he):(1'h0)] wire197;
  reg [(4'hf):(1'h0)] reg81 = (1'h0);
  reg [(4'he):(1'h0)] reg80 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg79 = (1'h0);
  reg [(2'h3):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg77 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar76 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg75 = (1'h0);
  reg [(4'hb):(1'h0)] reg74 = (1'h0);
  reg [(4'hf):(1'h0)] reg73 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar72 = (1'h0);
  reg [(5'h10):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar70 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg69 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar68 = (1'h0);
  reg [(5'h11):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg66 = (1'h0);
  reg [(5'h10):(1'h0)] reg65 = (1'h0);
  reg signed [(4'he):(1'h0)] reg64 = (1'h0);
  reg [(4'hf):(1'h0)] forvar63 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg62 = (1'h0);
  reg [(4'hc):(1'h0)] reg61 = (1'h0);
  reg [(3'h5):(1'h0)] reg60 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire59;
  wire [(4'hd):(1'h0)] wire57;
  wire signed [(5'h10):(1'h0)] wire28;
  wire [(5'h13):(1'h0)] wire27;
  wire [(5'h10):(1'h0)] wire410;
  wire [(5'h11):(1'h0)] wire563;
  wire [(5'h13):(1'h0)] wire569;
  wire signed [(4'ha):(1'h0)] wire570;
  assign y = {reg667,
                 forvar659,
                 reg658,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 forvar658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 forvar651,
                 reg650,
                 reg649,
                 reg648,
                 forvar647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 forvar642,
                 reg641,
                 forvar640,
                 wire639,
                 reg638,
                 reg637,
                 forvar636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 forvar630,
                 reg629,
                 reg628,
                 reg627,
                 forvar626,
                 reg625,
                 forvar624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 forvar618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 forvar612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 forvar605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 forvar599,
                 forvar598,
                 wire597,
                 reg596,
                 reg595,
                 reg594,
                 forvar593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 forvar587,
                 reg586,
                 forvar585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg577,
                 reg576,
                 forvar575,
                 reg574,
                 reg573,
                 wire572,
                 wire567,
                 wire566,
                 wire565,
                 wire561,
                 wire197,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 forvar76,
                 reg75,
                 reg74,
                 reg73,
                 forvar72,
                 reg71,
                 forvar70,
                 reg63,
                 reg69,
                 forvar68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 forvar63,
                 reg62,
                 reg61,
                 reg60,
                 wire59,
                 wire57,
                 wire28,
                 wire27,
                 wire410,
                 wire563,
                 wire569,
                 wire570,
                 (1'h0)};
  assign wire27 = wire23[(4'ha):(3'h5)];
  assign wire28 = (($unsigned((wire23 ^~ wire24)) ?
                          $signed((wire26[(3'h7):(3'h7)] == (wire27 >> wire24))) : ((8'ha4) ^ $unsigned(wire27))) ?
                      $unsigned(wire27[(1'h1):(1'h0)]) : wire25[(3'h7):(3'h5)]);
  module29 modinst58 (wire57, clk, wire23, wire27, wire26, wire28);
  assign wire59 = ($signed((~^$unsigned($unsigned(wire25)))) ?
                      wire24[(1'h0):(1'h0)] : wire24[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg60 <= ($signed(wire27) ? wire57 : wire25);
      reg61 = wire28;
      reg62 = (~|((8'ha3) >> ((wire26 ?
          (wire57 * wire24) : wire57) >>> $signed($unsigned(wire57)))));
      if (wire57[(4'hc):(3'h7)])
        begin
          for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
            begin
              reg64 <= (7'h44);
              reg65 <= ($signed(wire25) < wire25);
              reg66 <= $unsigned((^~reg60));
              reg67 = (({wire59[(1'h0):(1'h0)]} ?
                  $signed($signed($unsigned((7'h42)))) : forvar63) | ((8'hbe) >>> (reg62[(2'h3):(1'h1)] - $signed((reg61 <<< (7'h41))))));
            end
          for (forvar68 = (1'h0); (forvar68 < (2'h2)); forvar68 = (forvar68 + (1'h1)))
            begin
              reg69 <= (!(-reg61[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          reg63 = (|(~&forvar63));
          if ({$signed(reg65),
              $unsigned({{reg65[(2'h2):(1'h1)]}, (&$unsigned((8'haf)))})})
            begin
              reg64 <= (wire57[(4'h8):(3'h7)] ?
                  forvar63[(1'h0):(1'h0)] : wire57);
              reg65 = wire24;
              reg66 = $signed($signed((reg62[(3'h4):(1'h0)] == wire28)));
            end
          else
            begin
              reg64 = $unsigned($unsigned($signed((forvar63[(3'h4):(2'h2)] != $signed(forvar63)))));
              reg65 <= ((~wire59) ?
                  (8'ha3) : (|("BefQbxKYquXCnM" ?
                      $signed($signed((8'hb0))) : ($signed(reg67) ?
                          forvar68 : $unsigned(reg63)))));
              reg66 = ((8'hba) ?
                  wire25 : ((^~(^~(!reg69))) | (~|$unsigned((~|reg65)))));
              reg67 <= ($signed(reg65) <= reg62);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar70 = (1'h0); (forvar70 < (2'h3)); forvar70 = (forvar70 + (1'h1)))
        begin
          reg71 <= ($unsigned($signed((|((8'h9c) ?
              reg64 : (8'hb8))))) <= $unsigned((reg62[(1'h0):(1'h0)] >= ((~^forvar68) ~^ (!(7'h40))))));
          for (forvar72 = (1'h0); (forvar72 < (2'h2)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 <= (^~(((reg62[(2'h2):(1'h0)] || (reg71 << forvar72)) ?
                      $signed((wire59 ?
                          wire28 : forvar70)) : wire25[(4'hf):(2'h3)]) ?
                  $signed(((+reg67) > reg61)) : $signed((forvar72 ?
                      (reg71 < forvar70) : $unsigned(reg71)))));
              reg74 <= reg69[(1'h0):(1'h0)];
              reg75 = reg60;
            end
          for (forvar76 = (1'h0); (forvar76 < (1'h1)); forvar76 = (forvar76 + (1'h1)))
            begin
              reg77 = ((+$signed(((^(8'ha7)) ?
                  {wire28,
                      reg61} : forvar70))) ^ {{$unsigned((reg65 ^~ reg66))},
                  reg74});
              reg78 <= ($signed(wire27[(2'h3):(1'h1)]) ?
                  ((8'hb1) ? reg66 : wire23) : ({{$unsigned((8'ha7))},
                          wire27[(1'h1):(1'h1)]} ?
                      $unsigned($signed((forvar72 ?
                          forvar68 : wire28))) : {$unsigned(""),
                          ((wire59 || forvar63) ^ $signed(reg61))}));
              reg79 = wire23[(5'h12):(1'h1)];
              reg80 = (^forvar70);
              reg81 = wire25;
            end
        end
    end
  module82 modinst198 (.y(wire197), .wire84(forvar68), .clk(clk), .wire83(reg81), .wire87(reg73), .wire85(reg77), .wire86(wire23));
  module199 modinst411 (wire410, clk, wire26, reg66, reg67, reg65, reg74);
  module412 modinst562 (wire561, clk, reg65, forvar76, reg63, wire27, reg81);
  module82 modinst564 (wire563, clk, reg64, reg61, reg71, wire27, reg65);
  assign wire565 = forvar72;
  assign wire566 = (8'hb6);
  module82 modinst568 (wire567, clk, wire197, wire27, reg73, reg80, reg75);
  assign wire569 = reg80[(4'h8):(1'h1)];
  module412 modinst571 (.wire417(reg74), .wire416(reg67), .clk(clk), .wire413(reg69), .wire415(reg80), .y(wire570), .wire414(wire566));
  assign wire572 = $signed($unsigned((~|$signed($unsigned(reg75)))));
  always
    @(posedge clk) begin
      reg573 <= reg73[(4'h8):(1'h1)];
      reg574 = wire572;
    end
  always
    @(posedge clk) begin
      for (forvar575 = (1'h0); (forvar575 < (3'h4)); forvar575 = (forvar575 + (1'h1)))
        begin
          reg576 <= (8'hbb);
          reg577 <= ((-reg61[(2'h3):(2'h2)]) ?
              wire28 : $unsigned($unsigned((-(~|wire410)))));
          reg578 <= reg63[(4'h9):(3'h4)];
          for (forvar579 = (1'h0); (forvar579 < (2'h3)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 <= (|(&{(~^reg80),
                  ((+forvar70) ? wire26[(4'hc):(2'h2)] : wire26)}));
              reg581 <= $unsigned((wire25 ?
                  reg66[(3'h7):(2'h2)] : reg577[(1'h0):(1'h0)]));
              reg582 = (wire569[(4'hd):(4'ha)] < (!"Bs22GU8z5wdRBWeQ"));
              reg583 <= wire28;
              reg584 <= (^~(^~("y1UxK7nPzBy6RRoYBab6" && $unsigned(reg62))));
            end
        end
      for (forvar585 = (1'h0); (forvar585 < (3'h4)); forvar585 = (forvar585 + (1'h1)))
        begin
          reg586 <= $signed(wire25);
          for (forvar587 = (1'h0); (forvar587 < (1'h1)); forvar587 = (forvar587 + (1'h1)))
            begin
              reg588 = {wire26, (~&$unsigned((-(reg73 ? reg61 : reg586))))};
              reg589 <= wire566;
              reg590 <= {((reg65 ?
                          $unsigned($unsigned(reg71)) : (forvar63[(2'h2):(1'h0)] ?
                              (&reg81) : {wire59, wire561})) ?
                      (~(~(!reg62))) : wire567[(2'h3):(1'h0)]),
                  ($signed($unsigned(reg64[(2'h3):(2'h2)])) ?
                      (reg69[(4'hc):(2'h3)] == (~&$signed(reg80))) : (((reg73 << reg79) ?
                          $unsigned(reg67) : (-(8'ha2))) < $signed({(8'ha7),
                          wire23})))};
              reg591 <= reg79;
            end
          reg592 <= (~($signed({reg71[(5'h10):(4'hc)],
              $unsigned(wire25)}) ^~ $signed((&$signed(wire567)))));
          for (forvar593 = (1'h0); (forvar593 < (3'h4)); forvar593 = (forvar593 + (1'h1)))
            begin
              reg594 <= ((wire570 ?
                  wire25[(4'he):(3'h4)] : $signed($unsigned((reg79 && reg573)))) > $unsigned(reg81));
            end
          reg595 = (forvar68[(3'h6):(1'h0)] ?
              wire570[(4'h8):(1'h0)] : ((reg589 ?
                      ($signed(reg81) ?
                          $unsigned((8'hbd)) : reg576[(2'h3):(2'h2)]) : ($signed(reg586) ?
                          (reg61 ? reg75 : reg588) : reg73)) ?
                  wire26[(4'ha):(1'h0)] : ($signed($unsigned(wire570)) <= $signed({reg592,
                      wire572}))));
        end
      reg596 <= (((((wire24 ? reg592 : reg62) ? $signed(wire24) : reg583) ?
          ((reg74 - forvar579) ?
              (reg588 < wire572) : (reg591 ?
                  reg590 : reg61)) : {forvar68[(4'ha):(1'h1)]}) <= (~(8'hb3))) || (((7'h41) ?
              $unsigned($signed((8'hbb))) : {wire197[(2'h2):(2'h2)]}) ?
          (reg66[(3'h5):(1'h0)] == {$signed(reg74)}) : ($unsigned(reg578) != reg60[(3'h4):(2'h3)])));
    end
  assign wire597 = reg66[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar598 = (1'h0); (forvar598 < (2'h2)); forvar598 = (forvar598 + (1'h1)))
        begin
          for (forvar599 = (1'h0); (forvar599 < (2'h3)); forvar599 = (forvar599 + (1'h1)))
            begin
              reg600 <= $signed(({(~|(wire569 == wire572)),
                      forvar575[(4'hd):(3'h5)]} ?
                  $unsigned((^$signed((8'h9e)))) : wire28[(5'h10):(4'he)]));
              reg601 = wire572;
              reg602 = (8'hb0);
              reg603 <= $unsigned({{reg576[(4'h8):(1'h0)],
                      (reg71 ? $signed((8'ha4)) : (reg600 - reg74))}});
              reg604 = $signed(wire28[(4'ha):(4'ha)]);
            end
          for (forvar605 = (1'h0); (forvar605 < (1'h1)); forvar605 = (forvar605 + (1'h1)))
            begin
              reg606 <= wire57[(2'h2):(2'h2)];
              reg607 = $unsigned($signed(forvar68[(4'ha):(1'h0)]));
              reg608 <= $signed((wire59 < (((!reg582) ?
                  (reg578 ?
                      reg73 : forvar585) : $signed(reg77)) | (forvar599 - (~&reg79)))));
              reg609 <= $signed($unsigned(reg80[(4'h8):(1'h0)]));
              reg610 = reg69;
            end
          reg611 <= (&reg595[(1'h1):(1'h0)]);
          for (forvar612 = (1'h0); (forvar612 < (1'h0)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 = "EC9WE3m3v2";
              reg614 <= (^reg78[(1'h0):(1'h0)]);
              reg615 <= $signed($unsigned({{(~forvar575)},
                  ((~|forvar68) != reg576)}));
              reg616 <= $unsigned(reg608[(1'h1):(1'h0)]);
              reg617 <= (|{((+(reg75 >>> wire570)) ^ $signed(wire410[(1'h0):(1'h0)])),
                  (~&({wire197} ? "EpulJpyf5AEeF" : $signed((8'ha9))))});
            end
          for (forvar618 = (1'h0); (forvar618 < (3'h4)); forvar618 = (forvar618 + (1'h1)))
            begin
              reg619 <= reg79[(2'h2):(1'h0)];
              reg620 <= $unsigned(reg616[(1'h1):(1'h0)]);
              reg621 = reg74[(3'h7):(2'h2)];
              reg622 = forvar68[(3'h5):(1'h1)];
              reg623 <= $signed($signed(wire565[(2'h3):(1'h0)]));
            end
        end
      for (forvar624 = (1'h0); (forvar624 < (2'h2)); forvar624 = (forvar624 + (1'h1)))
        begin
          reg625 <= (((((reg573 ? reg78 : wire27) ^ "C7ZM7qgFJGd") ?
                  reg71 : $signed({(7'h44), reg622})) & $signed(reg66)) ?
              (forvar598 + $signed((reg60[(1'h0):(1'h0)] <= {reg574,
                  wire566}))) : $unsigned("vwihMdZkiTo"));
          for (forvar626 = (1'h0); (forvar626 < (2'h2)); forvar626 = (forvar626 + (1'h1)))
            begin
              reg627 = (("IA2qetRpwPMrXVlax" <<< ((^$unsigned(forvar579)) >= ((reg78 == reg81) ?
                      (~^reg591) : {(8'haf)}))) ?
                  $signed((wire566 ?
                      (~&(|reg608)) : (8'hbf))) : (reg589 << $unsigned(reg614[(3'h6):(1'h0)])));
              reg628 <= $unsigned(forvar612);
              reg629 <= (^"x4lRwzOpzGm");
            end
          for (forvar630 = (1'h0); (forvar630 < (1'h1)); forvar630 = (forvar630 + (1'h1)))
            begin
              reg631 = ((wire597 ?
                      {$unsigned(reg629[(4'hd):(3'h4)])} : "VfXz") ?
                  (~^wire23[(4'h8):(2'h2)]) : $unsigned((~^((reg80 ?
                          wire410 : (8'hb5)) ?
                      (&forvar63) : $signed((8'hbe))))));
              reg632 <= $signed(forvar605);
              reg633 <= $unsigned((({(8'ha2), {wire567}} + ((forvar624 ?
                      (7'h42) : (8'ha3)) ~^ $unsigned(wire23))) ?
                  $unsigned(wire25) : (+$unsigned(wire28[(4'hf):(4'hc)]))));
              reg634 <= (8'h9e);
              reg635 <= ({(^wire24), ($signed((~reg616)) <= {reg595})} ?
                  wire597[(4'hc):(2'h3)] : (~^$unsigned($signed($signed(reg621)))));
            end
          for (forvar636 = (1'h0); (forvar636 < (2'h3)); forvar636 = (forvar636 + (1'h1)))
            begin
              reg637 <= $signed((reg62[(2'h2):(1'h1)] - "bpaWuPEadVis"));
            end
        end
      reg638 = ({$signed($unsigned({forvar636}))} + wire565);
    end
  assign wire639 = (~&(&(|(reg613 ? (reg588 * reg74) : $unsigned(reg628)))));
  always
    @(posedge clk) begin
      for (forvar640 = (1'h0); (forvar640 < (1'h0)); forvar640 = (forvar640 + (1'h1)))
        begin
          reg641 = (8'hb3);
        end
      for (forvar642 = (1'h0); (forvar642 < (3'h4)); forvar642 = (forvar642 + (1'h1)))
        begin
          if ($signed(forvar624))
            begin
              reg643 <= reg584[(2'h3):(2'h3)];
              reg644 <= $unsigned(reg614);
              reg645 <= reg66[(1'h0):(1'h0)];
              reg646 <= (reg634 >>> reg582);
            end
          else
            begin
              reg643 <= {((8'ha1) == reg584[(3'h5):(2'h2)]),
                  reg582[(2'h2):(2'h2)]};
              reg644 <= reg586;
              reg645 <= reg601[(1'h1):(1'h1)];
              reg646 <= ("15l16AST" ?
                  "FPGEc" : ((8'ha8) ?
                      ({(forvar618 | reg602)} ?
                          (wire24 ?
                              $unsigned(reg75) : (reg603 ?
                                  reg625 : reg77)) : forvar587) : ("B3OMzh0OFTL3Tp" < ((~&reg589) ?
                          $signed(reg81) : reg592))));
            end
          for (forvar647 = (1'h0); (forvar647 < (3'h4)); forvar647 = (forvar647 + (1'h1)))
            begin
              reg648 = "a1J";
              reg649 <= (reg625 >>> (8'hb1));
              reg650 <= (~|(8'hb0));
            end
          for (forvar651 = (1'h0); (forvar651 < (1'h1)); forvar651 = (forvar651 + (1'h1)))
            begin
              reg652 = $signed($unsigned($signed($unsigned((!reg600)))));
              reg653 = $signed($signed(reg61[(3'h6):(3'h4)]));
              reg654 <= $signed($signed(((~&(~^reg590)) - ((reg620 - reg577) ?
                  $unsigned(reg71) : wire567))));
              reg655 <= (-reg583);
              reg656 <= {($signed({(reg63 ?
                          forvar579 : forvar647)}) | $unsigned({(reg582 ?
                          reg649 : (8'hbe))}))};
            end
          reg657 <= ($signed((reg62[(3'h4):(2'h3)] >= (((7'h43) * (8'haf)) || reg607))) ?
              $unsigned((reg615[(4'ha):(1'h1)] ~^ $unsigned($unsigned(reg649)))) : reg641);
        end
      if ($signed(reg582))
        begin
          for (forvar658 = (1'h0); (forvar658 < (2'h3)); forvar658 = (forvar658 + (1'h1)))
            begin
              reg659 <= (-$unsigned({$unsigned(forvar605[(3'h6):(1'h0)])}));
              reg660 <= ("" ? (7'h43) : (wire23 ^ (^(~$signed(reg632)))));
              reg661 <= {(+((reg637[(2'h3):(1'h0)] <= forvar612) ?
                      (&((7'h40) && forvar605)) : forvar599[(1'h0):(1'h0)]))};
            end
          reg662 <= ({reg615[(4'hc):(2'h2)]} ^~ $unsigned(reg615));
          if ($signed($unsigned((|reg80))))
            begin
              reg663 <= (((|{(forvar599 ? reg81 : reg632),
                      ((8'hb1) * reg589)}) >>> ((reg623 < $signed(wire565)) ?
                      {reg589,
                          reg69[(4'ha):(3'h4)]} : ($unsigned(forvar70) <<< reg62[(1'h1):(1'h0)]))) ?
                  "O69YFOHWn0Z9hyNvqLp" : wire572[(3'h6):(1'h1)]);
              reg664 = reg577[(1'h1):(1'h1)];
              reg665 = wire570[(3'h4):(1'h1)];
              reg666 <= (($unsigned((reg75[(3'h7):(1'h1)] + $signed(reg614))) ?
                      $unsigned(($unsigned(wire24) || (reg608 <= wire569))) : $signed(((!wire565) ?
                          wire27 : $signed(reg580)))) ?
                  ($signed((~^$signed(reg623))) * $unsigned((reg625 ?
                      "ozolu" : $unsigned(reg596)))) : reg590[(1'h0):(1'h0)]);
            end
          else
            begin
              reg663 <= (~(~&reg616[(4'h8):(2'h2)]));
            end
        end
      else
        begin
          reg658 <= ($unsigned(wire567) ?
              $unsigned((reg606[(2'h2):(1'h0)] ?
                  (~&(wire569 ? reg638 : (8'hab))) : ($signed(reg632) ?
                      wire26 : reg635))) : ((forvar72[(1'h0):(1'h0)] ?
                  forvar579 : ((forvar618 <= reg634) - $unsigned((8'ha7)))) > forvar624[(5'h14):(5'h10)]));
          for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= $unsigned($signed((reg80 ? reg653 : (~^(!forvar575)))));
            end
        end
      reg667 <= (7'h42);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module412
#( parameter param559 = ((((((8'hb9) ? (8'hba) : (8'ha7)) ? {(8'ha8), (7'h44)} : (&(8'ha5))) ? {((8'h9f) ? (8'hb7) : (8'h9d)), (^~(8'hb1))} : ((~^(8'h9d)) ? (^~(8'hb3)) : (^(7'h43)))) + (&(~|((8'ha9) ? (8'hb7) : (8'hb8))))) <<< ((-((8'ha8) <= {(8'hb9)})) ? (~&(+((8'ha6) ? (7'h42) : (8'h9c)))) : (~|(((8'hbc) ? (8'hb0) : (8'hbf)) ? ((8'ha5) ? (8'h9f) : (8'hbe)) : (-(8'hb8))))))
, parameter param560 = (~|((param559 ? (param559 ? {param559} : (param559 ? param559 : param559)) : ((param559 || (8'hab)) >>> (~|param559))) - (&(param559 ? param559 : param559)))) )
(y, clk, wire417, wire416, wire415, wire414, wire413);
  output wire [(32'h665):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire417;
  input wire [(4'he):(1'h0)] wire416;
  input wire signed [(3'h7):(1'h0)] wire415;
  input wire [(5'h13):(1'h0)] wire414;
  input wire [(4'hc):(1'h0)] wire413;
  wire signed [(3'h6):(1'h0)] wire558;
  wire signed [(3'h7):(1'h0)] wire557;
  wire signed [(3'h5):(1'h0)] wire556;
  reg signed [(4'hc):(1'h0)] reg555 = (1'h0);
  reg [(4'ha):(1'h0)] reg554 = (1'h0);
  reg signed [(4'he):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg552 = (1'h0);
  reg [(5'h13):(1'h0)] forvar551 = (1'h0);
  reg [(3'h4):(1'h0)] reg550 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg549 = (1'h0);
  reg [(4'he):(1'h0)] reg548 = (1'h0);
  reg [(5'h14):(1'h0)] reg547 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg546 = (1'h0);
  reg [(3'h7):(1'h0)] forvar545 = (1'h0);
  wire [(5'h10):(1'h0)] wire544;
  wire [(4'ha):(1'h0)] wire543;
  reg [(5'h14):(1'h0)] reg542 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg541 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar540 = (1'h0);
  reg [(4'hc):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg538 = (1'h0);
  reg [(4'hb):(1'h0)] reg537 = (1'h0);
  reg [(3'h7):(1'h0)] reg536 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar535 = (1'h0);
  reg [(5'h10):(1'h0)] reg534 = (1'h0);
  reg [(4'ha):(1'h0)] reg533 = (1'h0);
  reg [(4'hf):(1'h0)] reg532 = (1'h0);
  reg [(4'hd):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg530 = (1'h0);
  reg [(2'h2):(1'h0)] reg527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg524 = (1'h0);
  reg [(5'h15):(1'h0)] reg529 = (1'h0);
  reg [(4'h9):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar527 = (1'h0);
  reg [(5'h12):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg525 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar524 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg523 = (1'h0);
  reg [(5'h13):(1'h0)] reg522 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire521;
  wire signed [(5'h15):(1'h0)] wire520;
  reg signed [(4'hc):(1'h0)] reg519 = (1'h0);
  reg [(3'h4):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar517 = (1'h0);
  reg [(4'h8):(1'h0)] reg516 = (1'h0);
  reg [(3'h6):(1'h0)] reg515 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg514 = (1'h0);
  reg [(5'h11):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg512 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar511 = (1'h0);
  reg [(3'h6):(1'h0)] reg510 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg509 = (1'h0);
  reg [(4'ha):(1'h0)] forvar508 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg507 = (1'h0);
  reg [(4'ha):(1'h0)] reg506 = (1'h0);
  reg [(3'h4):(1'h0)] reg505 = (1'h0);
  reg [(4'h8):(1'h0)] reg504 = (1'h0);
  reg [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(5'h11):(1'h0)] reg502 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar501 = (1'h0);
  reg [(3'h6):(1'h0)] reg500 = (1'h0);
  reg [(4'hb):(1'h0)] reg499 = (1'h0);
  reg [(4'hd):(1'h0)] reg498 = (1'h0);
  reg [(4'hb):(1'h0)] reg497 = (1'h0);
  reg [(4'hf):(1'h0)] reg496 = (1'h0);
  reg signed [(4'he):(1'h0)] reg495 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg494 = (1'h0);
  reg [(5'h13):(1'h0)] reg493 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg492 = (1'h0);
  reg [(4'hc):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar490 = (1'h0);
  reg [(3'h4):(1'h0)] reg489 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg488 = (1'h0);
  reg [(3'h4):(1'h0)] forvar487 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar486 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg484 = (1'h0);
  reg [(4'hf):(1'h0)] reg483 = (1'h0);
  reg [(4'hb):(1'h0)] reg482 = (1'h0);
  reg [(4'hc):(1'h0)] reg481 = (1'h0);
  reg [(4'ha):(1'h0)] forvar480 = (1'h0);
  reg [(4'h9):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg478 = (1'h0);
  reg [(4'hb):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg476 = (1'h0);
  reg [(5'h12):(1'h0)] forvar475 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar474 = (1'h0);
  reg [(3'h5):(1'h0)] reg456 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg472 = (1'h0);
  reg [(4'hb):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg470 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar468 = (1'h0);
  reg [(3'h7):(1'h0)] reg467 = (1'h0);
  reg [(4'hd):(1'h0)] reg466 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg463 = (1'h0);
  reg [(4'h8):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg460 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg457 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar456 = (1'h0);
  reg signed [(4'he):(1'h0)] reg455 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg454 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar451 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg450 = (1'h0);
  reg [(3'h6):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar448 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg447 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg446 = (1'h0);
  reg [(2'h3):(1'h0)] forvar445 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg444 = (1'h0);
  reg [(5'h11):(1'h0)] reg443 = (1'h0);
  reg [(5'h10):(1'h0)] reg442 = (1'h0);
  reg [(4'h9):(1'h0)] forvar441 = (1'h0);
  reg [(4'h9):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg435 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg434 = (1'h0);
  reg [(5'h11):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg432 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg431 = (1'h0);
  reg [(4'hd):(1'h0)] reg430 = (1'h0);
  reg [(4'ha):(1'h0)] forvar429 = (1'h0);
  reg [(5'h11):(1'h0)] reg428 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg427 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar426 = (1'h0);
  reg [(4'h9):(1'h0)] reg419 = (1'h0);
  reg [(2'h2):(1'h0)] reg425 = (1'h0);
  reg [(3'h5):(1'h0)] reg424 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg423 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg422 = (1'h0);
  reg [(4'ha):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg420 = (1'h0);
  reg [(4'ha):(1'h0)] forvar419 = (1'h0);
  wire [(4'ha):(1'h0)] wire418;
  assign y = {wire558,
                 wire557,
                 wire556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 forvar551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 forvar545,
                 wire544,
                 wire543,
                 reg542,
                 reg541,
                 forvar540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 forvar535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg527,
                 reg524,
                 reg529,
                 reg528,
                 forvar527,
                 reg526,
                 reg525,
                 forvar524,
                 reg523,
                 reg522,
                 wire521,
                 wire520,
                 reg519,
                 reg518,
                 forvar517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 forvar511,
                 reg510,
                 reg509,
                 forvar508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 forvar490,
                 reg489,
                 reg488,
                 forvar487,
                 forvar486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 forvar475,
                 forvar474,
                 reg456,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 forvar468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 forvar456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 forvar451,
                 reg450,
                 reg449,
                 forvar448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 reg443,
                 reg442,
                 forvar441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 forvar429,
                 reg428,
                 reg427,
                 forvar426,
                 reg419,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 forvar419,
                 wire418,
                 (1'h0)};
  assign wire418 = wire417;
  always
    @(posedge clk) begin
      if ({$unsigned(($unsigned("TZr8THSPh0Hezokq3S4") ~^ wire417[(4'h8):(3'h7)]))})
        begin
          for (forvar419 = (1'h0); (forvar419 < (2'h3)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 = ($signed({wire413[(3'h6):(1'h0)],
                      ($unsigned((8'hb1)) ?
                          wire416[(1'h1):(1'h0)] : (forvar419 - wire413))}) ?
                  ({(-$unsigned(forvar419)), $unsigned({wire413})} ?
                      (|((forvar419 ^~ wire416) >> (8'ha0))) : (+(|wire415[(3'h5):(2'h2)]))) : wire417[(4'ha):(4'ha)]);
              reg421 = (^reg420);
              reg422 = $signed((|reg420));
              reg423 = $unsigned((wire418 ? reg422[(4'hc):(4'hc)] : reg420));
            end
          reg424 = {$signed((((wire416 ?
                  forvar419 : wire418) ^ $signed(reg422)) >>> $unsigned(wire413)))};
          reg425 = (((((wire413 - wire414) ?
                      reg420[(2'h2):(1'h0)] : $unsigned(reg420)) ?
                  wire415 : forvar419) == wire415[(2'h2):(1'h0)]) ?
              (8'hbf) : {$unsigned((8'ha2)),
                  (((reg420 <= reg421) ?
                          (reg424 ?
                              wire417 : wire416) : forvar419[(4'h8):(3'h6)]) ?
                      (reg424 * (!reg421)) : forvar419[(2'h2):(1'h1)])});
        end
      else
        begin
          reg419 = $unsigned($unsigned(($unsigned($unsigned(reg421)) ~^ (reg421[(2'h3):(1'h1)] ?
              (forvar419 >> wire417) : (^~reg423)))));
        end
      for (forvar426 = (1'h0); (forvar426 < (2'h2)); forvar426 = (forvar426 + (1'h1)))
        begin
          reg427 <= $unsigned({$signed($signed(reg424[(2'h2):(2'h2)]))});
          reg428 = ((wire417 ?
              "QoCm" : (~(~&(reg420 ?
                  wire413 : reg423)))) | (((wire415[(3'h6):(3'h6)] == (wire418 <<< wire416)) ?
                  (((8'ha7) ? reg425 : wire413) ?
                      (reg420 ?
                          (7'h43) : reg422) : $signed(wire415)) : forvar419[(3'h4):(2'h3)]) ?
              ({(&forvar426), (reg424 ? forvar419 : reg421)} ?
                  ("zB8ZStm" ?
                      "LDA7gbTbOFuG76tM" : (~(8'haf))) : {reg423[(3'h6):(1'h1)]}) : ((|(8'hbf)) ^ ((wire413 ?
                      wire415 : (8'hb9)) ?
                  wire418 : (^~wire415)))));
          for (forvar429 = (1'h0); (forvar429 < (3'h4)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 <= $unsigned((((reg420[(4'h9):(3'h7)] >>> (reg428 ?
                  wire416 : wire418)) < $unsigned($unsigned(forvar429))) < {((8'hac) ?
                      (-reg420) : reg423[(3'h4):(1'h0)])}));
              reg431 = (~$unsigned(((~|$unsigned(wire418)) * wire413[(1'h0):(1'h0)])));
              reg432 = {$unsigned(reg422)};
              reg433 <= wire415[(3'h7):(2'h3)];
            end
          if ("8OnK")
            begin
              reg434 = ((reg428[(4'h9):(4'h8)] ?
                      $unsigned((wire416 == (reg419 ?
                          reg423 : wire416))) : forvar429[(3'h4):(1'h1)]) ?
                  "6spHvTw" : "AcSvlmtMoudg9");
              reg435 = $unsigned(wire413[(1'h1):(1'h1)]);
              reg436 <= (~|$unsigned(reg432[(2'h2):(1'h0)]));
              reg437 <= $signed((^(-wire418)));
              reg438 = wire417[(3'h5):(2'h2)];
            end
          else
            begin
              reg434 <= (((wire418 < $unsigned($unsigned(reg437))) ~^ (wire415[(3'h7):(1'h0)] ?
                      reg424 : $unsigned(reg431))) ?
                  {$signed(({reg434, (8'hb8)} | (^~reg421))),
                      reg427[(3'h7):(3'h7)]} : $unsigned(($signed($signed(reg422)) >> reg419[(3'h5):(1'h1)])));
              reg435 <= (8'hba);
              reg436 <= $signed((8'ha5));
              reg437 <= wire414;
              reg438 <= (reg422[(2'h3):(2'h3)] ? reg425 : "OoSFnIbbKOE");
            end
        end
      reg439 = ((reg427[(2'h2):(1'h0)] >>> reg435) ?
          (!{$unsigned($signed((8'h9f)))}) : ($unsigned(($unsigned((8'hb2)) ~^ (reg423 - reg422))) ?
              wire413 : (wire413[(4'ha):(2'h2)] > $signed(reg420))));
      reg440 = $unsigned((((-$unsigned(wire417)) ?
          reg428 : (+(~&reg433))) << ($signed($signed(wire416)) ?
          ({forvar426, (8'ha4)} ?
              (+reg421) : $signed(wire413)) : $unsigned($signed((8'ha8))))));
    end
  always
    @(posedge clk) begin
      for (forvar441 = (1'h0); (forvar441 < (1'h0)); forvar441 = (forvar441 + (1'h1)))
        begin
          reg442 <= (wire415 >= wire417);
          reg443 <= (&reg430);
          reg444 <= reg422;
          for (forvar445 = (1'h0); (forvar445 < (1'h0)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= reg424;
            end
          reg447 = reg446[(2'h3):(1'h1)];
        end
      for (forvar448 = (1'h0); (forvar448 < (2'h2)); forvar448 = (forvar448 + (1'h1)))
        begin
          reg449 = (&({reg443[(4'hc):(4'h9)]} ?
              $signed((forvar448 ? reg436 : reg438[(1'h1):(1'h1)])) : reg437));
          reg450 <= $unsigned($signed((reg419[(2'h2):(2'h2)] * $unsigned($unsigned(forvar419)))));
          for (forvar451 = (1'h0); (forvar451 < (1'h1)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 <= (reg427[(3'h4):(2'h3)] << $unsigned($unsigned(reg430)));
            end
          reg453 = $unsigned(($unsigned(wire416) | (($signed(reg440) ^~ (wire417 | reg437)) ?
              $signed(forvar451) : wire416)));
          if ("UpoAuQtGyA2lf7")
            begin
              reg454 <= reg432;
              reg455 <= ((($unsigned((reg434 ?
                      reg420 : reg431)) << {reg444[(3'h4):(1'h1)]}) != $signed($signed(reg431[(2'h2):(1'h1)]))) ?
                  (8'ha5) : $signed({$signed(reg447[(3'h4):(1'h0)])}));
            end
          else
            begin
              reg454 = (~^(reg423[(4'ha):(1'h1)] ?
                  $signed(((~^(7'h40)) | (reg455 ~^ reg449))) : ("0ERcD0fw97TA2d" >>> $unsigned(((8'hab) ?
                      reg453 : reg436)))));
            end
        end
      if (((~^$signed(((~reg442) >> (8'had)))) ?
          (7'h43) : (($signed($unsigned(wire414)) ?
                  reg428 : (reg436[(4'h8):(2'h2)] >>> (^~reg422))) ?
              {$unsigned(reg431[(1'h0):(1'h0)]),
                  (((8'hac) && forvar441) + (forvar419 ?
                      (8'ha8) : (8'ha4)))} : $signed($unsigned((^~reg436))))))
        begin
          for (forvar456 = (1'h0); (forvar456 < (3'h4)); forvar456 = (forvar456 + (1'h1)))
            begin
              reg457 <= (^~("l1CPeayhuNnKA" & $signed((reg447[(1'h0):(1'h0)] ?
                  ((7'h44) ? (7'h42) : reg453) : (~|reg447)))));
              reg458 = $signed($signed($unsigned($unsigned(reg431[(1'h0):(1'h0)]))));
              reg459 <= (({"maOxiXS0VAVAy4Y"} ?
                  (~$signed($signed(reg435))) : reg424) && $unsigned(wire417[(4'hb):(3'h5)]));
              reg460 = (^~((reg455[(3'h4):(1'h0)] ?
                      $signed($unsigned(reg427)) : ((~&reg424) ?
                          (reg457 ? reg425 : reg435) : reg420[(2'h3):(2'h3)])) ?
                  (~|{(wire414 ? reg455 : reg419),
                      (reg443 * forvar419)}) : ($unsigned((reg442 ?
                      reg455 : reg443)) + reg428)));
            end
          reg461 <= (!wire414);
          reg462 <= (($signed({$unsigned(wire414), reg428}) ?
                  $signed({$unsigned(reg430), $unsigned(wire415)}) : reg421) ?
              wire416[(4'h9):(2'h2)] : (~^forvar451[(2'h3):(2'h3)]));
          if ($signed((^~$unsigned(wire414))))
            begin
              reg463 <= $unsigned(reg427[(1'h0):(1'h0)]);
              reg464 = (^~(^~(((~reg420) - $signed(reg444)) >= ((reg461 ^~ reg460) ?
                  $signed(reg427) : forvar448))));
              reg465 = ($unsigned($unsigned($signed((~^reg459)))) == $unsigned($unsigned($unsigned(((8'hb0) <= wire413)))));
              reg466 = reg454[(1'h0):(1'h0)];
              reg467 <= $unsigned((-$signed($unsigned((reg438 >>> reg455)))));
            end
          else
            begin
              reg463 <= reg463;
              reg464 <= $signed(forvar451[(2'h2):(1'h1)]);
              reg465 <= ($unsigned("uW68") > reg447);
            end
          for (forvar468 = (1'h0); (forvar468 < (2'h3)); forvar468 = (forvar468 + (1'h1)))
            begin
              reg469 = reg460;
              reg470 = $signed(reg458);
              reg471 <= {$signed({reg457})};
              reg472 = $signed((+$signed($unsigned(reg453))));
              reg473 <= $unsigned({(reg470[(1'h1):(1'h1)] && forvar429[(2'h2):(1'h0)])});
            end
        end
      else
        begin
          reg456 = (~^reg422);
        end
    end
  always
    @(posedge clk) begin
      for (forvar474 = (1'h0); (forvar474 < (3'h4)); forvar474 = (forvar474 + (1'h1)))
        begin
          for (forvar475 = (1'h0); (forvar475 < (2'h3)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 = ((~reg419) | (^(8'ha4)));
              reg477 = $signed({$signed(wire415[(2'h3):(2'h2)])});
            end
          reg478 = $signed(reg456);
          if ((-reg443[(4'h8):(2'h2)]))
            begin
              reg479 = $unsigned(reg470[(3'h6):(2'h2)]);
            end
          else
            begin
              reg479 = $signed($unsigned((((8'hbb) ?
                      $unsigned(reg433) : reg479[(1'h0):(1'h0)]) ?
                  reg452[(3'h7):(2'h2)] : $signed($signed(reg427)))));
            end
          for (forvar480 = (1'h0); (forvar480 < (3'h4)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= forvar480;
              reg482 <= reg479[(4'h9):(1'h0)];
              reg483 = reg447[(3'h7):(3'h4)];
              reg484 <= wire415[(1'h0):(1'h0)];
              reg485 <= {forvar468[(4'he):(4'he)]};
            end
        end
      for (forvar486 = (1'h0); (forvar486 < (3'h4)); forvar486 = (forvar486 + (1'h1)))
        begin
          for (forvar487 = (1'h0); (forvar487 < (1'h1)); forvar487 = (forvar487 + (1'h1)))
            begin
              reg488 = {(~$unsigned(reg484)), forvar445[(2'h2):(2'h2)]};
              reg489 <= reg477;
            end
          for (forvar490 = (1'h0); (forvar490 < (2'h2)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 <= {$unsigned((reg485 ? (7'h43) : reg470)),
                  $signed($unsigned($signed((reg439 | wire418))))};
              reg492 <= $unsigned((reg466[(3'h5):(2'h3)] <= ($unsigned(reg438[(1'h1):(1'h1)]) ?
                  $signed((7'h42)) : reg470)));
              reg493 <= forvar480;
              reg494 = ($signed((8'h9f)) ~^ $unsigned(forvar480));
              reg495 <= $signed((reg446[(4'h8):(1'h1)] ?
                  $signed(reg430) : reg478[(4'he):(4'ha)]));
            end
          if ((reg454 << $signed($unsigned($unsigned((~|reg461))))))
            begin
              reg496 <= ($unsigned(($unsigned($signed(forvar474)) ?
                  $unsigned((reg423 ?
                      (8'ha1) : reg424)) : ((~^reg422) ~^ (reg494 > reg470)))) >> (reg471 ?
                  ((reg476[(4'hd):(4'hc)] < {reg473}) >> ($signed(forvar456) ^~ reg462[(4'h8):(3'h6)])) : (+(8'hac))));
              reg497 = (({$signed($signed(reg421)),
                      (8'ha9)} & $unsigned({(reg435 && reg454)})) ?
                  ((+$unsigned((forvar475 <= reg496))) ?
                      $unsigned(reg436) : (~&$unsigned($signed((8'hae))))) : forvar445[(2'h2):(1'h1)]);
              reg498 <= $unsigned($unsigned(reg463));
              reg499 <= {(+(((reg432 << reg484) & (reg473 ?
                          forvar441 : reg424)) ?
                      (^(reg433 == reg482)) : $unsigned(reg450))),
                  {$signed($signed(reg473)), ($signed((7'h44)) * reg472)}};
              reg500 = $unsigned((($unsigned("GfhcGEf") ?
                  "cT66wrRqq2gKmua" : reg439) ^ {reg478}));
            end
          else
            begin
              reg496 <= reg438[(1'h1):(1'h1)];
              reg497 = (-{(reg495[(4'h9):(2'h3)] >>> reg455),
                  (((reg447 >= reg431) ?
                      (|reg428) : $unsigned(reg461)) < $unsigned($signed((7'h42))))});
              reg498 <= (^~reg478);
              reg499 = $signed(wire416);
            end
          for (forvar501 = (1'h0); (forvar501 < (2'h3)); forvar501 = (forvar501 + (1'h1)))
            begin
              reg502 = reg488;
              reg503 = ({$signed((+reg427[(2'h3):(2'h3)]))} - $unsigned(reg449));
              reg504 = {{"yMOLQB"}, {(^~reg446[(2'h3):(1'h1)])}};
            end
          reg505 <= (reg493[(3'h6):(2'h2)] ?
              $signed((^~(reg456[(2'h2):(2'h2)] ^~ (reg476 ?
                  reg498 : reg458)))) : reg422[(4'hf):(3'h4)]);
        end
      reg506 = (~(($signed((forvar451 >>> forvar451)) ?
              (|reg483[(4'h8):(3'h7)]) : reg466) ?
          {$signed((8'hbf))} : {reg456, (~|reg505)}));
      reg507 <= {((reg452 ?
                  $signed((reg496 >>> reg504)) : ($signed(reg458) < (reg423 ?
                      reg472 : (8'hae)))) ?
              "W3M2u" : $unsigned((&(~reg458)))),
          ($unsigned(reg442[(4'hb):(4'ha)]) <= $signed($signed((~&(8'ha8)))))};
      for (forvar508 = (1'h0); (forvar508 < (1'h1)); forvar508 = (forvar508 + (1'h1)))
        begin
          if (((~^($unsigned(reg495) >= reg447[(3'h6):(1'h0)])) | forvar419[(3'h6):(3'h6)]))
            begin
              reg509 = ((-(-(reg453 ? $signed((8'hb5)) : {reg473, reg422}))) ?
                  ($unsigned($signed((~&reg479))) ?
                      (~&reg450[(3'h6):(1'h1)]) : (((forvar426 ?
                              wire416 : reg457) <= reg497) ?
                          ($signed(reg457) ?
                              (reg472 >>> reg443) : (forvar490 ~^ reg439)) : reg450[(3'h6):(3'h6)])) : (8'hbd));
            end
          else
            begin
              reg509 <= (forvar448 >> (forvar441 >> reg482[(4'h8):(3'h6)]));
              reg510 <= (&reg464);
            end
          for (forvar511 = (1'h0); (forvar511 < (2'h2)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 = {((|forvar468[(4'hb):(1'h0)]) >>> (reg439 ?
                      forvar501[(4'h9):(3'h6)] : $signed((reg427 <<< reg450)))),
                  reg465};
              reg513 <= (((-reg424) ? forvar508[(2'h2):(1'h0)] : (8'hb6)) ?
                  "s" : forvar474[(3'h5):(1'h0)]);
              reg514 <= $unsigned((^~(reg453 ?
                  (^~{reg507}) : $signed(reg421))));
              reg515 <= (^~$signed((reg488[(3'h6):(3'h4)] ?
                  (reg510 || (forvar451 ? reg457 : reg469)) : (reg495 ?
                      $unsigned(reg484) : $unsigned(reg493)))));
              reg516 = ((+(!$signed(wire418[(3'h7):(3'h4)]))) >>> $signed($signed(reg500)));
            end
          for (forvar517 = (1'h0); (forvar517 < (2'h3)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 <= (^(&forvar474));
              reg519 <= (+$signed(reg446[(4'h9):(3'h6)]));
            end
        end
    end
  assign wire520 = $signed($signed($signed("v")));
  assign wire521 = ({(~|$signed((forvar441 <= (8'hb3)))),
                           {(+(wire520 - reg515))}} ?
                       "iPl5SbsHZ" : $signed(((~|(~&forvar448)) | $signed($unsigned((8'hb6))))));
  always
    @(posedge clk) begin
      if (($signed(($signed(reg461) && $unsigned((reg516 ?
              forvar501 : reg420)))) ?
          forvar508[(3'h7):(3'h4)] : (forvar490 ?
              (~|(~(-reg515))) : $signed(forvar501))))
        begin
          reg522 = ((|$unsigned(($unsigned(reg433) ~^ (8'hb2)))) << (~$signed($signed(((8'ha8) == (8'ha9))))));
          reg523 = (+(^~$signed({$unsigned(reg492)})));
          for (forvar524 = (1'h0); (forvar524 < (1'h1)); forvar524 = (forvar524 + (1'h1)))
            begin
              reg525 = $signed($unsigned(wire414[(5'h11):(4'ha)]));
            end
          reg526 <= $unsigned(reg424[(3'h4):(3'h4)]);
          for (forvar527 = (1'h0); (forvar527 < (1'h0)); forvar527 = (forvar527 + (1'h1)))
            begin
              reg528 <= $unsigned((($unsigned($signed(reg498)) ?
                      $unsigned({(7'h41), reg507}) : (forvar475 ?
                          "V4LdK8FoFDm9" : (!reg463))) ?
                  (~reg481) : forvar448));
              reg529 <= reg430[(2'h2):(2'h2)];
            end
        end
      else
        begin
          reg522 = ((forvar419 > (+reg453[(3'h5):(2'h2)])) ^ (~|($unsigned(reg483) != (reg428[(4'hc):(3'h6)] | {(7'h44),
              (8'hbf)}))));
          if (($signed((^~$signed(reg491[(3'h6):(2'h3)]))) ?
              (($unsigned($signed(reg489)) ?
                      reg420[(4'h9):(3'h7)] : $unsigned(forvar451)) ?
                  "J6wWwWp96" : $signed($signed($unsigned((8'ha9))))) : ("7Puas01deE8E3" ?
                  {reg500[(3'h5):(2'h3)],
                      $unsigned($signed(reg512))} : $signed("o6YeBAFHe8aBZK6aYv"))))
            begin
              reg523 = (&forvar426[(3'h4):(2'h3)]);
              reg524 = {reg502, reg497};
              reg525 <= {((^($unsigned((8'h9c)) ?
                      $signed(reg470) : (reg507 ?
                          reg462 : reg465))) | (^reg438[(2'h2):(1'h0)])),
                  (((~^$signed(reg419)) ?
                      ((forvar474 != reg434) ?
                          reg507[(1'h1):(1'h0)] : (!(7'h40))) : $unsigned($unsigned(wire417))) + (-$signed(reg481)))};
              reg526 = ((!$signed(((~|reg433) | (^(8'ha5))))) | (-(!$signed($unsigned(reg496)))));
            end
          else
            begin
              reg523 = $unsigned(reg422);
              reg524 = $unsigned({(8'h9e),
                  $unsigned((&((8'hbe) ? wire521 : reg489)))});
            end
          if ((~&($unsigned("EO2QnlK00Kn4OD4NKOhW") ?
              ((+reg454[(2'h2):(2'h2)]) ?
                  (+$signed(forvar468)) : ($unsigned(reg453) ?
                      ((8'hbb) ^~ reg461) : reg478)) : ((+(reg478 - forvar419)) ?
                  $unsigned(forvar456) : {(reg494 ? (8'hb0) : (8'ha3)),
                      $unsigned((8'ha4))}))))
            begin
              reg527 <= {"ucmWzZ42T", reg442[(4'he):(4'hd)]};
            end
          else
            begin
              reg527 <= (^$unsigned((reg482[(2'h3):(2'h2)] + wire413[(4'hb):(4'h8)])));
              reg528 = (!forvar474[(2'h3):(2'h3)]);
              reg529 <= $unsigned({($unsigned((&reg450)) || reg479[(1'h0):(1'h0)])});
            end
          if ($signed((({(reg453 + reg478),
              (~(8'hb0))} * "YF6YxvRy6thG") + $unsigned($signed({forvar486,
              reg484})))))
            begin
              reg530 = (^reg440[(1'h1):(1'h0)]);
              reg531 = $unsigned({$unsigned(((+reg476) <= $signed(reg485))),
                  (&forvar480[(3'h6):(1'h0)])});
              reg532 = (|reg450);
              reg533 = reg460;
              reg534 = ((((-(reg522 ?
                          forvar429 : reg485)) || ($unsigned((8'hb2)) * (wire417 ?
                          reg500 : reg462))) ?
                      $signed((8'ha1)) : reg516) ?
                  $unsigned((forvar429[(4'h9):(3'h6)] | ($signed((8'hb9)) ?
                      (forvar511 ?
                          reg459 : reg454) : reg449[(3'h4):(1'h0)]))) : ((8'hb4) + (reg471 ?
                      ({reg497,
                          reg526} & reg446[(4'h8):(3'h7)]) : $unsigned((!wire416)))));
            end
          else
            begin
              reg530 = {(~{((reg515 ^~ reg446) > "fw7GfQ4dr55J"),
                      (!(~&reg419))}),
                  reg516};
              reg531 <= ($unsigned((-reg498)) ?
                  ((-((&(8'hab)) >>> reg512[(3'h5):(3'h5)])) >= $unsigned((~^$signed(reg505)))) : ((~&reg433) || (reg515[(2'h3):(2'h2)] + $signed($signed(reg497)))));
              reg532 = (|(8'ha8));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar535 = (1'h0); (forvar535 < (3'h4)); forvar535 = (forvar535 + (1'h1)))
        begin
          if (reg435[(1'h1):(1'h0)])
            begin
              reg536 <= ($signed((-$signed((reg425 ? forvar419 : reg503)))) ?
                  $signed((reg478[(3'h7):(3'h5)] & reg469[(4'h9):(1'h0)])) : ($unsigned(forvar445[(2'h2):(1'h1)]) >> reg489));
            end
          else
            begin
              reg536 <= $unsigned((+reg464));
              reg537 <= (|(!$unsigned(reg456)));
            end
          reg538 <= $unsigned($signed(($unsigned(reg478[(3'h5):(2'h3)]) >>> reg422)));
        end
      reg539 <= reg505;
      for (forvar540 = (1'h0); (forvar540 < (2'h3)); forvar540 = (forvar540 + (1'h1)))
        begin
          reg541 = $signed($unsigned((8'ha3)));
          if ({(reg502[(4'hd):(4'h9)] ?
                  $signed(($signed(forvar468) ?
                      $signed(reg537) : {forvar448})) : $unsigned((((8'h9d) ?
                      reg485 : (8'hb9)) << $unsigned((8'hb3)))))})
            begin
              reg542 <= (~((-(!reg450[(3'h5):(3'h4)])) ?
                  (+("" ^ $signed(reg534))) : (8'ha1)));
            end
          else
            begin
              reg542 <= forvar475;
            end
        end
    end
  assign wire543 = reg427;
  assign wire544 = (-$unsigned($unsigned(((reg458 ?
                       reg519 : reg440) ~^ (~&reg484)))));
  always
    @(posedge clk) begin
      for (forvar545 = (1'h0); (forvar545 < (2'h3)); forvar545 = (forvar545 + (1'h1)))
        begin
          if (reg539)
            begin
              reg546 <= $unsigned(((+reg518) < reg499[(1'h0):(1'h0)]));
              reg547 = $signed($unsigned(reg421[(3'h6):(3'h5)]));
              reg548 <= ($signed($unsigned(reg533[(1'h1):(1'h0)])) == reg497);
              reg549 <= ($unsigned((^reg476[(3'h4):(2'h3)])) ^ (+(~|"F7Si")));
            end
          else
            begin
              reg546 = reg471[(3'h5):(3'h4)];
              reg547 <= reg504;
              reg548 = (reg433 ?
                  (^reg548) : (reg548 ?
                      (~forvar426) : {{{(8'hb5)}}, $signed({forvar445})}));
              reg549 = (reg541 << ({{reg473}, reg458} >> $unsigned(((forvar511 ?
                      reg432 : reg537) ?
                  (reg423 >= (8'ha5)) : $signed(wire543)))));
              reg550 = $signed((~|((&reg463) ?
                  (8'hae) : forvar511[(4'h9):(2'h2)])));
            end
          for (forvar551 = (1'h0); (forvar551 < (2'h3)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 <= $signed((7'h43));
              reg553 <= (-reg444);
              reg554 = $unsigned(({{(forvar490 - reg529), reg424}} ?
                  $unsigned(reg456[(1'h0):(1'h0)]) : reg538));
              reg555 <= (~reg529[(5'h14):(3'h4)]);
            end
        end
    end
  assign wire556 = (-$signed("BRKmUhdKQiSH"));
  assign wire557 = {forvar501};
  assign wire558 = reg424[(3'h5):(3'h4)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module199
#( parameter param409 = (((~&(8'hb5)) ? (7'h41) : {(-((7'h44) ? (8'hbf) : (8'ha5)))}) ? (((((8'ha8) ? (7'h42) : (8'hb5)) ? (~^(8'ha8)) : (~(8'ha7))) ? {(~&(8'hbe)), ((8'hb1) ? (8'h9d) : (8'h9c))} : ((&(8'haf)) | ((8'hbf) || (8'ha6)))) ? (((-(8'hb3)) ? {(7'h44)} : (8'ha1)) ? (((8'hbf) < (8'hbf)) ? ((8'hb8) ? (8'ha6) : (8'hb3)) : (~(7'h44))) : (~^((8'hac) << (7'h40)))) : ((+((7'h43) & (8'hb4))) >= (^~((8'ha4) ? (8'h9e) : (8'hab))))) : {(~^(((8'h9e) > (8'hbb)) - ((8'h9d) ? (8'hb6) : (8'hb7))))}) )
(y, clk, wire204, wire203, wire202, wire201, wire200);
  output wire [(32'h978):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire204;
  input wire signed [(3'h7):(1'h0)] wire203;
  input wire [(5'h11):(1'h0)] wire202;
  input wire signed [(5'h10):(1'h0)] wire201;
  input wire [(3'h4):(1'h0)] wire200;
  wire signed [(3'h5):(1'h0)] wire408;
  reg signed [(2'h2):(1'h0)] reg407 = (1'h0);
  reg [(5'h12):(1'h0)] reg406 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg404 = (1'h0);
  reg [(5'h12):(1'h0)] reg403 = (1'h0);
  reg [(5'h10):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg401 = (1'h0);
  reg [(4'hc):(1'h0)] reg400 = (1'h0);
  reg [(4'hd):(1'h0)] reg399 = (1'h0);
  reg [(4'h9):(1'h0)] reg398 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg397 = (1'h0);
  reg [(4'hc):(1'h0)] reg396 = (1'h0);
  reg [(5'h14):(1'h0)] reg395 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg388 = (1'h0);
  reg [(3'h7):(1'h0)] forvar386 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg383 = (1'h0);
  reg [(4'hb):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg393 = (1'h0);
  reg [(2'h2):(1'h0)] reg392 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg389 = (1'h0);
  reg [(4'h8):(1'h0)] forvar388 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg387 = (1'h0);
  reg [(4'hf):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg385 = (1'h0);
  reg [(5'h10):(1'h0)] reg384 = (1'h0);
  reg [(3'h6):(1'h0)] forvar383 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg382 = (1'h0);
  reg [(3'h6):(1'h0)] reg381 = (1'h0);
  reg [(3'h6):(1'h0)] reg380 = (1'h0);
  wire [(4'hf):(1'h0)] wire379;
  reg signed [(5'h14):(1'h0)] reg378 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg376 = (1'h0);
  reg [(4'hd):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg374 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar373 = (1'h0);
  reg [(4'hc):(1'h0)] reg372 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar371 = (1'h0);
  reg [(4'h8):(1'h0)] reg370 = (1'h0);
  reg [(5'h12):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg368 = (1'h0);
  reg [(5'h11):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar366 = (1'h0);
  reg [(5'h15):(1'h0)] forvar365 = (1'h0);
  wire [(2'h2):(1'h0)] wire364;
  wire [(3'h5):(1'h0)] wire363;
  wire signed [(4'hc):(1'h0)] wire362;
  reg signed [(2'h2):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar360 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg359 = (1'h0);
  reg [(4'hf):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg356 = (1'h0);
  reg [(3'h6):(1'h0)] reg355 = (1'h0);
  reg [(2'h3):(1'h0)] forvar354 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg352 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar351 = (1'h0);
  reg [(4'h8):(1'h0)] reg350 = (1'h0);
  reg [(4'hb):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar347 = (1'h0);
  reg [(4'hc):(1'h0)] reg346 = (1'h0);
  reg [(4'ha):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg343 = (1'h0);
  reg [(3'h4):(1'h0)] reg342 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg341 = (1'h0);
  reg [(5'h12):(1'h0)] forvar340 = (1'h0);
  reg [(3'h6):(1'h0)] reg340 = (1'h0);
  reg [(2'h2):(1'h0)] reg339 = (1'h0);
  reg [(3'h5):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg337 = (1'h0);
  reg [(3'h4):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg335 = (1'h0);
  reg [(4'ha):(1'h0)] reg334 = (1'h0);
  wire signed [(4'he):(1'h0)] wire333;
  wire [(2'h3):(1'h0)] wire332;
  reg signed [(5'h11):(1'h0)] reg331 = (1'h0);
  reg [(3'h4):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg329 = (1'h0);
  reg [(4'hf):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg327 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar326 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg325 = (1'h0);
  reg [(4'hc):(1'h0)] reg324 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg323 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar322 = (1'h0);
  reg [(4'h8):(1'h0)] reg321 = (1'h0);
  reg [(5'h11):(1'h0)] reg320 = (1'h0);
  reg [(4'h9):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg315 = (1'h0);
  reg [(5'h14):(1'h0)] forvar314 = (1'h0);
  reg [(2'h2):(1'h0)] reg313 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg311 = (1'h0);
  reg [(3'h6):(1'h0)] forvar310 = (1'h0);
  reg [(5'h15):(1'h0)] forvar309 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg307 = (1'h0);
  reg [(5'h10):(1'h0)] reg294 = (1'h0);
  reg [(4'h9):(1'h0)] reg306 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg303 = (1'h0);
  reg [(3'h5):(1'h0)] reg302 = (1'h0);
  reg [(5'h11):(1'h0)] reg301 = (1'h0);
  reg [(4'he):(1'h0)] reg300 = (1'h0);
  reg [(4'hb):(1'h0)] reg299 = (1'h0);
  reg [(4'h9):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg297 = (1'h0);
  reg [(5'h10):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg295 = (1'h0);
  reg [(5'h13):(1'h0)] forvar294 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg293 = (1'h0);
  reg [(5'h11):(1'h0)] reg292 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg291 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg289 = (1'h0);
  reg [(4'h8):(1'h0)] forvar288 = (1'h0);
  reg [(5'h15):(1'h0)] reg287 = (1'h0);
  reg [(5'h13):(1'h0)] reg286 = (1'h0);
  reg [(5'h13):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] forvar284 = (1'h0);
  reg [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg282 = (1'h0);
  reg signed [(4'he):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar280 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg279 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg277 = (1'h0);
  reg [(2'h2):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar274 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg273 = (1'h0);
  reg [(5'h12):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar269 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg268 = (1'h0);
  reg [(4'h8):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg263 = (1'h0);
  reg [(4'h9):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar261 = (1'h0);
  reg [(4'h9):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar259 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(4'h8):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar253 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg252 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg251 = (1'h0);
  reg [(4'hc):(1'h0)] reg250 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg249 = (1'h0);
  reg [(3'h4):(1'h0)] reg248 = (1'h0);
  reg [(5'h14):(1'h0)] forvar247 = (1'h0);
  reg [(4'hb):(1'h0)] reg246 = (1'h0);
  reg [(4'hc):(1'h0)] reg245 = (1'h0);
  reg [(5'h10):(1'h0)] reg244 = (1'h0);
  reg [(4'h8):(1'h0)] reg243 = (1'h0);
  reg [(3'h7):(1'h0)] forvar242 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar241 = (1'h0);
  wire [(4'he):(1'h0)] wire240;
  wire signed [(4'hd):(1'h0)] wire239;
  wire signed [(4'hc):(1'h0)] wire238;
  reg [(2'h2):(1'h0)] reg237 = (1'h0);
  reg [(4'hc):(1'h0)] reg236 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg235 = (1'h0);
  reg [(3'h7):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar233 = (1'h0);
  reg [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg231 = (1'h0);
  reg [(3'h5):(1'h0)] forvar230 = (1'h0);
  reg [(5'h12):(1'h0)] forvar229 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg228 = (1'h0);
  reg [(4'hc):(1'h0)] reg227 = (1'h0);
  reg [(4'hd):(1'h0)] forvar226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg223 = (1'h0);
  reg [(3'h5):(1'h0)] reg222 = (1'h0);
  reg [(4'h8):(1'h0)] forvar221 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar220 = (1'h0);
  reg [(5'h12):(1'h0)] reg219 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg215 = (1'h0);
  reg [(5'h10):(1'h0)] reg214 = (1'h0);
  reg [(2'h2):(1'h0)] reg213 = (1'h0);
  reg [(2'h3):(1'h0)] reg212 = (1'h0);
  reg [(4'hf):(1'h0)] reg211 = (1'h0);
  reg [(2'h2):(1'h0)] reg210 = (1'h0);
  reg [(3'h6):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg208 = (1'h0);
  reg [(5'h10):(1'h0)] forvar207 = (1'h0);
  reg [(5'h15):(1'h0)] forvar206 = (1'h0);
  wire [(4'hd):(1'h0)] wire205;
  assign y = {wire408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg388,
                 forvar386,
                 reg383,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 forvar388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 forvar383,
                 reg382,
                 reg381,
                 reg380,
                 wire379,
                 reg378,
                 forvar377,
                 reg376,
                 reg375,
                 reg374,
                 forvar373,
                 reg372,
                 forvar371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 forvar366,
                 forvar365,
                 wire364,
                 wire363,
                 wire362,
                 reg361,
                 forvar360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 forvar354,
                 reg353,
                 reg352,
                 forvar351,
                 reg350,
                 reg349,
                 reg348,
                 forvar347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 forvar340,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 wire333,
                 wire332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 forvar326,
                 reg325,
                 reg324,
                 reg323,
                 forvar322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 reg317,
                 reg316,
                 reg315,
                 forvar314,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 forvar309,
                 reg308,
                 reg307,
                 reg294,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 forvar294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 forvar288,
                 reg287,
                 reg286,
                 reg285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 forvar280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 forvar274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 forvar269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 forvar261,
                 reg260,
                 forvar259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 forvar253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 forvar247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 forvar242,
                 forvar241,
                 wire240,
                 wire239,
                 wire238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 reg232,
                 reg231,
                 forvar230,
                 forvar229,
                 reg228,
                 reg227,
                 forvar226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 forvar221,
                 forvar220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 forvar207,
                 forvar206,
                 wire205,
                 (1'h0)};
  assign wire205 = wire203[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar206 = (1'h0); (forvar206 < (1'h0)); forvar206 = (forvar206 + (1'h1)))
        begin
          for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 = $signed(wire203[(3'h6):(1'h0)]);
              reg209 <= ((!{{(|wire200)},
                  ((-forvar206) ^ reg208[(4'h8):(3'h4)])}) || wire204);
              reg210 = forvar207;
              reg211 <= ((|wire205) ?
                  ((!(~(|reg208))) ?
                      $signed((~^wire203)) : {{wire201, (reg208 - (8'hb3))},
                          (~&$signed((8'hbe)))}) : ($unsigned((wire201[(4'ha):(3'h6)] <= (&(8'hbb)))) + (+$signed($signed(reg208)))));
              reg212 = wire204[(5'h10):(1'h1)];
            end
          reg213 <= {reg208[(2'h2):(1'h0)],
              (((+wire205) >> "iv1PKQP1t") ?
                  $unsigned($unsigned((&forvar207))) : $signed((^reg208)))};
          reg214 = (({(~(^~wire200)),
                      (wire205[(1'h0):(1'h0)] ^~ forvar206[(4'h9):(3'h5)])} ?
                  $signed((reg212 & (wire200 >>> reg212))) : $unsigned(wire204)) ?
              ($signed(wire201) ?
                  $signed($unsigned((~^reg213))) : (8'haf)) : wire201);
          if (wire202[(2'h2):(2'h2)])
            begin
              reg215 <= ((($unsigned(reg210) != (wire205[(4'hb):(2'h2)] ?
                      ((8'h9c) ?
                          wire203 : forvar206) : $signed(wire202))) >= $signed({(forvar207 < forvar207),
                      (^(8'ha0))})) ?
                  ({reg213} ?
                      ($signed(wire203) ?
                          $unsigned((wire204 ?
                              wire203 : forvar206)) : ($unsigned(wire203) >= (8'hb8))) : $signed({((8'ha9) + reg208)})) : $unsigned(({(reg211 ?
                          reg212 : forvar207),
                      {forvar207}} + {$unsigned(reg213),
                      wire202[(1'h1):(1'h1)]})));
              reg216 = ($signed((($unsigned(wire201) ?
                      $unsigned(reg208) : $signed(wire200)) - reg215[(1'h1):(1'h1)])) ?
                  reg213 : $signed(reg209));
              reg217 = ((8'hb5) ?
                  $unsigned(wire202) : ((+wire200[(2'h2):(1'h0)]) ?
                      wire205 : wire201[(3'h7):(3'h5)]));
              reg218 <= {{wire203}};
            end
          else
            begin
              reg215 = wire203;
              reg216 <= (^~((^~$unsigned((reg213 ? reg209 : reg208))) ?
                  reg214[(2'h2):(2'h2)] : (|$signed((8'had)))));
              reg217 <= $unsigned($unsigned({((^reg218) ?
                      {(8'ha2), forvar206} : reg210[(2'h2):(1'h0)])}));
            end
          reg219 <= (reg210[(2'h2):(1'h1)] ?
              $signed((reg209[(3'h6):(3'h5)] ?
                  $signed((reg218 ^~ reg212)) : "CwOGEagrTvyw9Ph4")) : (!((^~(wire201 > reg215)) ^ $signed($unsigned(wire202)))));
        end
      for (forvar220 = (1'h0); (forvar220 < (3'h4)); forvar220 = (forvar220 + (1'h1)))
        begin
          for (forvar221 = (1'h0); (forvar221 < (1'h0)); forvar221 = (forvar221 + (1'h1)))
            begin
              reg222 = reg217;
              reg223 <= $signed((reg219[(3'h5):(1'h0)] ?
                  reg215[(2'h2):(1'h0)] : reg215[(4'ha):(4'h9)]));
            end
          reg224 <= $unsigned($signed((~^(^(wire200 && wire200)))));
          reg225 <= reg213[(2'h2):(1'h1)];
        end
      for (forvar226 = (1'h0); (forvar226 < (2'h3)); forvar226 = (forvar226 + (1'h1)))
        begin
          reg227 = reg222[(1'h0):(1'h0)];
          reg228 <= reg219;
        end
      for (forvar229 = (1'h0); (forvar229 < (2'h2)); forvar229 = (forvar229 + (1'h1)))
        begin
          for (forvar230 = (1'h0); (forvar230 < (1'h1)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 <= wire201[(3'h6):(2'h3)];
            end
          reg232 <= $unsigned((^wire202));
          for (forvar233 = (1'h0); (forvar233 < (1'h1)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 = ({{$unsigned((reg215 ? reg217 : forvar221)),
                          $unsigned((reg228 <= reg219))}} ?
                  (($unsigned(reg222[(2'h3):(1'h0)]) ?
                          $unsigned($signed(reg228)) : "n6pfYGwzTq3s7XUH") ?
                      (^~$unsigned(reg210)) : forvar221[(1'h0):(1'h0)]) : forvar220);
              reg235 <= $signed(($signed("kB") ?
                  $unsigned(((reg216 << reg222) <= (~|(8'haa)))) : (8'h9c)));
            end
          reg236 <= "Zt7OocoM4hIO";
        end
      if (($unsigned((8'hbc)) ?
          (^reg234) : $signed({$unsigned($unsigned(forvar229)),
              forvar229[(4'ha):(1'h0)]})))
        begin
          reg237 = $signed((reg212 ?
              (~^(8'ha8)) : $unsigned((forvar229[(3'h6):(3'h6)] ^~ (forvar221 ?
                  reg209 : reg214)))));
        end
      else
        begin
          reg237 = ($unsigned(((wire203 && (reg216 - reg234)) ?
                  (8'hb5) : ((~^forvar206) ~^ $signed(reg223)))) ?
              $unsigned($unsigned(($signed(reg222) ?
                  "wRUtE0T" : (reg208 ?
                      reg237 : wire205)))) : ((!$signed(reg211[(4'he):(1'h0)])) ?
                  $unsigned(reg225) : $unsigned(((8'hb7) ?
                      {wire205} : (reg225 ? reg218 : reg236)))));
        end
    end
  assign wire238 = (~^({$unsigned($unsigned(forvar221)),
                           (+(wire203 ? reg210 : reg231))} ?
                       ($signed($signed(wire200)) ^ reg217[(4'hb):(1'h1)]) : reg227));
  assign wire239 = reg223[(5'h13):(4'h9)];
  assign wire240 = $signed((8'hbc));
  always
    @(posedge clk) begin
      for (forvar241 = (1'h0); (forvar241 < (1'h0)); forvar241 = (forvar241 + (1'h1)))
        begin
          for (forvar242 = (1'h0); (forvar242 < (3'h4)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 = (($unsigned((+$signed(reg214))) * $signed(reg227)) ?
                  (^~$unsigned(wire202)) : (&$signed("QXEVSKm")));
              reg244 = reg234[(1'h0):(1'h0)];
            end
        end
      if (forvar226)
        begin
          reg245 = reg214[(3'h7):(2'h2)];
        end
      else
        begin
          reg245 <= $signed((((~^(reg228 ? (8'h9e) : reg216)) ?
              $unsigned($unsigned(forvar230)) : $signed($signed(wire240))) ^~ $unsigned({wire200[(2'h3):(1'h0)]})));
          if (reg218[(4'ha):(1'h1)])
            begin
              reg246 = $unsigned(reg237);
            end
          else
            begin
              reg246 <= reg223[(4'hf):(4'h9)];
            end
          for (forvar247 = (1'h0); (forvar247 < (1'h0)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= $signed($signed($unsigned($signed({reg234}))));
              reg249 = reg222[(1'h0):(1'h0)];
              reg250 <= $unsigned((^~forvar221[(1'h0):(1'h0)]));
              reg251 <= $signed($unsigned((8'ha0)));
            end
          reg252 <= ($unsigned((((~^(7'h41)) >>> (reg249 >= reg243)) >> ((forvar220 <= reg225) > {reg224,
              wire240}))) >> forvar220);
        end
      if ({(($signed({reg251}) ?
              ((reg235 >>> wire202) ?
                  (forvar230 == reg234) : (8'hb1)) : forvar226) >> ($signed((^~forvar207)) ?
              reg210 : $unsigned($signed(reg210))))})
        begin
          for (forvar253 = (1'h0); (forvar253 < (1'h0)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= (^~{{reg213[(1'h0):(1'h0)],
                      {(reg218 ? reg246 : (8'hb3)), reg237}},
                  {$unsigned((|reg224))}});
              reg255 = $signed((-$signed($unsigned($signed((8'h9d))))));
              reg256 = (reg210[(1'h0):(1'h0)] ?
                  $signed((({(8'ha2), forvar230} ?
                          (~&reg209) : $signed(forvar233)) ?
                      (forvar242[(3'h7):(3'h4)] >= reg249[(4'h8):(1'h0)]) : ($unsigned(reg235) <<< "7BaHNNopwiI8m1KQQd"))) : (reg255 - forvar247));
            end
          reg257 <= (~reg250[(3'h7):(2'h3)]);
        end
      else
        begin
          for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= reg213[(1'h0):(1'h0)];
              reg255 <= reg237;
              reg256 = reg252[(3'h6):(2'h2)];
            end
          reg257 <= (^reg256[(2'h3):(1'h0)]);
          reg258 <= ($signed($signed(($unsigned(reg249) ?
              reg257[(4'hf):(3'h5)] : wire203[(3'h7):(1'h1)]))) | ((~^(~^forvar247)) && ({(reg223 && (7'h42)),
                  $signed(reg209)} ?
              reg213 : (!(forvar207 <= reg214)))));
          for (forvar259 = (1'h0); (forvar259 < (1'h1)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 = $unsigned({wire203});
            end
        end
      for (forvar261 = (1'h0); (forvar261 < (2'h2)); forvar261 = (forvar261 + (1'h1)))
        begin
          if (reg234)
            begin
              reg262 <= (|(reg235 <<< reg258[(1'h0):(1'h0)]));
            end
          else
            begin
              reg262 <= ($unsigned($signed(forvar241[(3'h6):(2'h3)])) - (~$signed((reg222[(1'h1):(1'h0)] - (forvar226 ~^ wire201)))));
              reg263 <= reg235[(5'h12):(3'h7)];
              reg264 <= (reg211[(2'h3):(2'h2)] ?
                  ($unsigned($unsigned(reg225)) <= (|forvar253[(3'h5):(1'h1)])) : (((+$unsigned(reg215)) ?
                          reg243[(3'h7):(3'h4)] : ({reg234, wire205} ?
                              (forvar242 ? reg217 : reg245) : {reg262,
                                  reg243})) ?
                      $unsigned(forvar226) : {{{reg219, reg232},
                              wire200[(3'h4):(3'h4)]}}));
              reg265 = reg219[(5'h10):(3'h7)];
              reg266 <= $signed($unsigned((-(^"YZyYiZh7I2zQ"))));
            end
          reg267 <= (+(^~reg223));
          reg268 <= $unsigned((-{({reg251} ? reg217[(4'hc):(3'h4)] : reg235)}));
          for (forvar269 = (1'h0); (forvar269 < (2'h2)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 <= $signed($signed({($signed(wire201) ?
                      (!reg267) : forvar253[(2'h3):(1'h1)])}));
              reg271 <= (("7m" ?
                  (~$signed($unsigned(reg248))) : $signed($signed({(8'hac)}))) * (~|({(reg236 ?
                          reg211 : reg210)} ?
                  reg222[(3'h5):(3'h4)] : $unsigned($unsigned((8'ha4))))));
              reg272 <= (forvar220[(2'h2):(2'h2)] ?
                  ($signed(((wire239 >= reg268) ? reg235 : wire239)) ?
                      $signed(reg252[(2'h3):(2'h3)]) : $signed($signed($signed(forvar242)))) : $signed(reg232[(2'h3):(1'h0)]));
              reg273 = $signed($unsigned($unsigned(((reg232 - (8'h9e)) ?
                  (forvar220 >= reg256) : ((8'ha9) ? reg250 : reg217)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg219[(4'hf):(3'h6)] | $signed({$signed((forvar247 > reg237))})))
        begin
          for (forvar274 = (1'h0); (forvar274 < (3'h4)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 <= ((8'haf) && $unsigned(reg228[(4'h9):(4'h9)]));
            end
          reg276 <= "s3s";
          reg277 <= (&($signed(((reg265 ? reg232 : (7'h40)) == (8'hb6))) ?
              wire200 : (^~$unsigned("l28"))));
        end
      else
        begin
          for (forvar274 = (1'h0); (forvar274 < (3'h4)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 = (((reg224 == ((reg214 ? wire239 : forvar220) ?
                          forvar247[(2'h3):(1'h0)] : wire203)) ?
                      $unsigned($unsigned((forvar242 ?
                          reg237 : forvar241))) : $signed(reg256)) ?
                  forvar229 : {reg272[(3'h4):(3'h4)]});
              reg276 = ($signed((((forvar259 <= reg250) ~^ (~^reg249)) != $unsigned($unsigned(forvar269)))) >> ((-(reg251[(1'h0):(1'h0)] <<< $signed((7'h41)))) >>> ($signed($unsigned((8'hb0))) > forvar261)));
              reg277 <= reg218;
            end
          if ("FaksNM77qmKzeK")
            begin
              reg278 = "Qa91Eq9QLv";
              reg279 = reg209;
            end
          else
            begin
              reg278 <= (($signed(reg218[(3'h4):(1'h1)]) ?
                  reg234 : (forvar242 >>> reg212[(2'h3):(2'h2)])) != ((8'hbb) ^~ $signed({reg244,
                  (wire203 <<< reg224)})));
              reg279 <= reg273[(4'h9):(3'h5)];
            end
          for (forvar280 = (1'h0); (forvar280 < (2'h3)); forvar280 = (forvar280 + (1'h1)))
            begin
              reg281 = $signed((($unsigned($signed(reg210)) >>> forvar261) ^~ $signed(forvar269[(4'hd):(4'h8)])));
              reg282 <= reg256;
              reg283 <= $signed({({{forvar274},
                      ((8'h9f) >>> reg282)} == (((7'h44) ?
                          forvar269 : (8'haf)) ?
                      {reg281, forvar253} : (reg249 ^~ reg214))),
                  (~&$unsigned($signed((7'h41))))});
            end
          for (forvar284 = (1'h0); (forvar284 < (3'h4)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 = forvar259[(4'hd):(4'h9)];
              reg286 <= $signed(reg252);
              reg287 <= {wire201,
                  ($signed($unsigned((reg236 ? reg282 : (8'hb3)))) ?
                      (8'hbe) : (reg243 ?
                          reg260 : (forvar241[(5'h12):(4'hb)] ?
                              wire201 : $signed(forvar233))))};
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
        begin
          if ($unsigned(((reg268[(3'h6):(3'h4)] || ($signed(reg244) ?
              (reg271 ?
                  reg215 : (8'h9c)) : reg244[(1'h1):(1'h1)])) != $signed({reg223[(5'h15):(1'h1)],
              ((8'hb8) ? reg258 : wire201)}))))
            begin
              reg289 <= (reg225[(1'h0):(1'h0)] ?
                  (reg248 ?
                      reg277[(1'h1):(1'h1)] : ($unsigned((forvar259 >>> (7'h42))) ?
                          (^$signed((8'hbf))) : ((wire238 ?
                                  reg215 : forvar284) ?
                              (&wire238) : (~&reg217)))) : ($unsigned((~(8'hbd))) ?
                      $signed(reg270) : (((+reg225) - $signed(reg273)) << $signed($unsigned(reg276)))));
              reg290 <= reg250;
              reg291 <= $signed(forvar274);
              reg292 <= (-$unsigned({(~|(~&reg254))}));
            end
          else
            begin
              reg289 <= $unsigned((&reg268));
              reg290 = "q";
            end
        end
      reg293 = $unsigned((reg285[(1'h0):(1'h0)] ?
          ((reg222 >>> (8'haf)) >>> $unsigned((reg260 && reg232))) : $unsigned((&(forvar241 ?
              (8'hbb) : forvar221)))));
    end
  always
    @(posedge clk) begin
      if ($unsigned("h"))
        begin
          for (forvar294 = (1'h0); (forvar294 < (3'h4)); forvar294 = (forvar294 + (1'h1)))
            begin
              reg295 <= reg291;
              reg296 <= ($signed($unsigned($unsigned((reg264 ?
                  forvar269 : reg237)))) != {($signed(wire202[(4'hb):(1'h0)]) ?
                      ((reg267 ?
                          (8'ha5) : reg273) ^~ $signed(forvar259)) : (~&reg268[(1'h1):(1'h0)])),
                  forvar288});
            end
          if (($signed(($signed(reg215[(2'h2):(1'h1)]) <<< ($unsigned((8'hbb)) ?
                  (wire240 > reg282) : {forvar284, reg235}))) ?
              reg222[(2'h3):(2'h2)] : (~&$signed(((forvar253 ?
                  reg236 : forvar280) & $unsigned(forvar247))))))
            begin
              reg297 <= $unsigned(reg281);
            end
          else
            begin
              reg297 <= $unsigned($signed((^~wire200[(1'h1):(1'h0)])));
              reg298 <= $signed(reg281);
              reg299 <= (((((reg212 ? reg211 : forvar280) ?
                          {(8'hab)} : (reg250 ? reg231 : reg292)) ?
                      ($unsigned(forvar229) ?
                          (8'hba) : $signed(reg213)) : reg296) == forvar274) ?
                  ($signed($unsigned($signed(wire239))) && reg216[(3'h5):(1'h0)]) : "b");
              reg300 <= ($unsigned((((|reg262) ?
                          (reg281 ^~ reg263) : (reg286 ? reg211 : reg222)) ?
                      (8'ha6) : reg235[(4'ha):(2'h2)])) ?
                  {forvar230} : reg272[(3'h7):(1'h0)]);
              reg301 <= reg275[(2'h2):(1'h1)];
            end
          if (($signed(forvar280) ?
              (&$unsigned((~&$signed(wire201)))) : (^~(&reg214[(4'h9):(1'h0)]))))
            begin
              reg302 <= (8'ha8);
              reg303 = $unsigned({(8'hb3),
                  ($signed((+reg275)) | $signed((~&reg271)))});
              reg304 = $unsigned(forvar269);
              reg305 <= $signed(forvar288[(3'h7):(1'h0)]);
              reg306 = (~^(-reg305[(3'h7):(3'h4)]));
            end
          else
            begin
              reg302 <= (|$unsigned((reg232[(1'h1):(1'h0)] ?
                  reg208[(4'hc):(3'h6)] : (~reg301))));
            end
        end
      else
        begin
          reg294 <= (({((reg224 ? reg272 : forvar269) <<< reg295),
                      "QgrWCBwb3dtqU9mZd4"} ?
                  reg256 : (~($signed(reg213) ?
                      (~|reg210) : $unsigned(forvar280)))) ?
              (&$signed($unsigned(wire200[(1'h1):(1'h0)]))) : (~|$signed($unsigned((~wire202)))));
          if ((((~^$unsigned($unsigned(reg278))) ?
              $unsigned({forvar220,
                  wire203[(3'h4):(1'h0)]}) : $unsigned(((reg222 ?
                      reg292 : (8'hac)) ?
                  (wire200 ?
                      reg257 : reg293) : (~reg249)))) == $unsigned(forvar207)))
            begin
              reg295 = forvar288[(3'h7):(2'h3)];
              reg296 <= ($unsigned(((|"sU6SwaAJs") & ($signed((8'h9d)) ?
                      (reg266 * forvar284) : $signed(wire239)))) ?
                  reg219 : $signed(((reg271 ?
                          $unsigned((8'ha5)) : $signed(reg235)) ?
                      (8'haa) : reg232)));
              reg297 = {$signed(($unsigned((reg235 ? (8'h9f) : forvar230)) ?
                      $signed({reg260,
                          reg303}) : ($unsigned(forvar242) >= (|reg213)))),
                  (reg306[(3'h6):(1'h0)] ?
                      (+{$unsigned(reg298),
                          reg277[(1'h1):(1'h1)]}) : $unsigned(($signed(reg212) ?
                          {reg237} : $signed(reg254))))};
              reg298 <= reg249;
            end
          else
            begin
              reg295 <= reg275[(4'h9):(2'h3)];
              reg296 <= reg236[(4'ha):(1'h0)];
              reg297 = (^~((reg296 ?
                  (8'hba) : {(reg210 ? reg292 : reg222),
                      forvar284}) ^ $unsigned(((reg277 << forvar269) ?
                  $unsigned(reg252) : reg296[(2'h3):(1'h0)]))));
            end
          reg299 = (($signed($signed(reg212)) ?
              (reg273 <= {reg215[(4'hb):(3'h6)]}) : forvar288) ^ $unsigned($unsigned(reg249)));
        end
      reg307 <= (~^{$unsigned(reg260), $signed(forvar206[(5'h14):(5'h13)])});
      reg308 = ((+(&{{reg295}, $signed(reg303)})) ?
          (~|reg296[(3'h7):(2'h3)]) : reg231);
      for (forvar309 = (1'h0); (forvar309 < (3'h4)); forvar309 = (forvar309 + (1'h1)))
        begin
          for (forvar310 = (1'h0); (forvar310 < (2'h3)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 <= ((~{reg285,
                  reg289[(3'h5):(3'h5)]}) && $signed((forvar220 ?
                  (^~$unsigned((8'hb5))) : $signed(reg299[(2'h3):(2'h2)]))));
              reg312 = ($unsigned(forvar247) <= $unsigned(forvar269[(4'hb):(4'hb)]));
              reg313 <= ($signed((!$signed(((8'ha3) >>> (8'ha4))))) & (~reg283));
            end
          for (forvar314 = (1'h0); (forvar314 < (1'h0)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg315 <= $unsigned(($unsigned({$unsigned(reg312)}) ?
                  $signed(((reg257 ? forvar226 : reg286) ?
                      $unsigned(reg265) : (reg308 ?
                          reg295 : (8'hb9)))) : (+$unsigned($unsigned((8'hb3))))));
              reg316 <= {reg249[(2'h2):(1'h1)],
                  ((^~(reg299 << (reg285 << reg213))) ?
                      $signed({(reg215 | reg265),
                          forvar288}) : (reg295 || {reg303,
                          $unsigned(reg237)}))};
              reg317 = reg307[(3'h7):(3'h6)];
            end
        end
      for (forvar318 = (1'h0); (forvar318 < (3'h4)); forvar318 = (forvar318 + (1'h1)))
        begin
          if ($unsigned((((|reg254[(1'h0):(1'h0)]) * reg317) && $signed({reg281[(4'hc):(4'ha)],
              reg218}))))
            begin
              reg319 <= (~|$signed($signed($signed($unsigned(reg211)))));
            end
          else
            begin
              reg319 = $signed($unsigned((~|({reg257} > $unsigned(forvar309)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg320 <= ((~^((wire238 ?
                  (reg260 ? reg218 : reg250) : (reg254 + forvar284)) ?
              reg218[(2'h3):(2'h3)] : ($unsigned(forvar314) ?
                  $signed((8'ha9)) : $signed(reg305)))) ?
          $signed(reg231[(5'h13):(4'hc)]) : wire203[(3'h6):(1'h1)]);
      reg321 <= (((reg245 ? reg210 : (reg290[(2'h3):(2'h3)] != "NNWI")) ?
          ({reg252[(1'h1):(1'h1)]} ?
              reg279 : reg266) : reg307[(4'hf):(4'hc)]) >= ($signed($signed((~^reg292))) & (!(forvar207 >> "PnmOGQqaUbXZrXkR"))));
      for (forvar322 = (1'h0); (forvar322 < (3'h4)); forvar322 = (forvar322 + (1'h1)))
        begin
          reg323 <= ({(8'h9c)} >> $unsigned(((~&$signed(reg308)) ?
              $unsigned(reg222[(3'h4):(2'h3)]) : $unsigned(reg298))));
          reg324 = {$signed(((&reg252) >= reg218)),
              ($unsigned(($signed(reg212) << reg258[(1'h1):(1'h0)])) ?
                  {({reg260, reg295} ?
                          (forvar322 ? reg228 : reg278) : {(8'ha1)}),
                      $unsigned(reg258)} : $signed((^~$unsigned(reg306))))};
          reg325 = (reg308[(3'h5):(1'h1)] * (^(-$unsigned((reg231 ?
              reg300 : (8'hb9))))));
          for (forvar326 = (1'h0); (forvar326 < (1'h0)); forvar326 = (forvar326 + (1'h1)))
            begin
              reg327 = reg210;
            end
          if ($signed((reg283[(2'h3):(1'h0)] ?
              $signed((~^(reg324 ^~ reg237))) : (~^reg273[(3'h5):(2'h2)]))))
            begin
              reg328 = forvar269;
              reg329 <= $unsigned((8'hb1));
              reg330 = (((-({reg264, reg210} << (forvar221 ?
                      forvar206 : reg275))) ?
                  (8'hb4) : (reg243[(3'h7):(3'h4)] <= (|reg295))) ^~ $signed((+(reg211[(1'h0):(1'h0)] ?
                  (reg299 ? reg287 : reg301) : ((8'ha9) ? wire205 : reg313)))));
              reg331 <= (^reg295);
            end
          else
            begin
              reg328 = $signed((~reg265));
              reg329 <= reg245;
              reg330 = $signed("JpmUtwpRYkfSvwJyt2i");
              reg331 = reg265;
            end
        end
    end
  assign wire332 = (reg278 ?
                       $unsigned(((~|forvar226) || $unsigned(reg294[(3'h6):(3'h4)]))) : ($unsigned((reg250 >>> (reg222 ?
                               (8'hb0) : (8'hb5)))) ?
                           ($unsigned((!reg294)) - $unsigned(reg214[(3'h4):(2'h2)])) : ($signed((reg315 * reg289)) || (&(^reg283)))));
  assign wire333 = $unsigned($signed((~|reg306)));
  always
    @(posedge clk) begin
      if (($unsigned($signed(($signed(forvar310) ?
              $unsigned((7'h44)) : {reg268}))) ?
          (|(~|($signed(reg300) == reg285))) : reg303[(3'h4):(2'h3)]))
        begin
          reg334 = ((forvar284 - "Qx0XiLXnxGf67") ?
              (reg211[(4'hf):(4'hb)] ?
                  (-reg287) : reg327) : $unsigned("HBR2bJd7Cewf7"));
        end
      else
        begin
          reg334 <= (~&$unsigned($signed(($unsigned(forvar314) * reg287[(2'h3):(1'h0)]))));
          if (forvar221)
            begin
              reg335 = (^($signed($unsigned($signed((8'hb1)))) ?
                  {({(8'hbe), forvar310} ? (~|forvar284) : $signed(reg297)),
                      reg256[(4'h8):(1'h0)]} : reg211[(3'h6):(3'h5)]));
            end
          else
            begin
              reg335 <= ((8'hb3) ?
                  $signed($signed($signed((!reg292)))) : $unsigned((!$signed(reg237[(1'h1):(1'h1)]))));
              reg336 <= (((({reg328} ?
                          ((8'ha2) - (8'hbd)) : $unsigned(wire200)) ?
                      reg279[(5'h14):(2'h3)] : reg254) << $unsigned(forvar207[(3'h4):(3'h4)])) ?
                  {$unsigned(((reg265 ? forvar242 : reg311) ?
                          $signed(forvar233) : {wire203, wire238})),
                      {forvar207[(4'hc):(2'h2)]}} : reg250);
              reg337 <= (~&(+reg311[(4'h9):(2'h2)]));
            end
          reg338 = reg266;
          reg339 = reg210;
        end
      if ($unsigned(reg323[(1'h0):(1'h0)]))
        begin
          reg340 <= ($signed((($signed(reg260) - $signed((8'hb5))) == reg324[(4'hc):(3'h5)])) != reg236[(3'h7):(2'h2)]);
        end
      else
        begin
          for (forvar340 = (1'h0); (forvar340 < (2'h2)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= reg317[(1'h1):(1'h1)];
            end
          if ($signed(($unsigned({(wire200 << reg340)}) >> (($signed(reg296) & (^(7'h41))) ?
              wire239 : (reg316[(1'h1):(1'h0)] ?
                  $unsigned(reg312) : (reg317 ? forvar253 : reg294))))))
            begin
              reg342 = reg296[(1'h1):(1'h1)];
              reg343 <= (8'hbb);
            end
          else
            begin
              reg342 = $unsigned(((~^(8'ha0)) < reg319[(3'h7):(1'h0)]));
              reg343 <= (|$unsigned($signed(reg330[(2'h2):(1'h0)])));
              reg344 <= (!($signed({forvar294[(5'h12):(4'ha)]}) ?
                  (((forvar314 ? wire239 : (8'hbb)) * (forvar242 ?
                      reg236 : reg319)) + ((reg256 ?
                      forvar288 : reg291) <<< {reg245})) : {reg251[(2'h2):(1'h0)]}));
              reg345 = {$unsigned(({reg248[(1'h0):(1'h0)]} ?
                      (&$unsigned(forvar253)) : reg330)),
                  (~^reg295)};
              reg346 <= $unsigned(wire200);
            end
          for (forvar347 = (1'h0); (forvar347 < (2'h3)); forvar347 = (forvar347 + (1'h1)))
            begin
              reg348 <= reg329;
              reg349 <= reg275;
              reg350 = "emEmvzahFqGmvoM1";
            end
        end
      for (forvar351 = (1'h0); (forvar351 < (1'h1)); forvar351 = (forvar351 + (1'h1)))
        begin
          reg352 <= reg294;
          reg353 <= (|reg312[(2'h3):(2'h2)]);
          for (forvar354 = (1'h0); (forvar354 < (3'h4)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 <= $unsigned($signed($signed({reg263[(2'h2):(1'h1)],
                  reg276})));
              reg356 <= (~|$signed(forvar226));
              reg357 = (~|reg350);
              reg358 <= {(-reg298[(3'h5):(1'h1)])};
            end
        end
      reg359 <= (~|reg323);
      for (forvar360 = (1'h0); (forvar360 < (3'h4)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 = ($unsigned({{$unsigned(wire332)}}) ^~ ((^~(~^reg319[(3'h6):(3'h6)])) ?
              ($signed($signed(forvar261)) <= (reg215[(4'h8):(3'h4)] ?
                  (!reg338) : reg248[(1'h0):(1'h0)])) : ((+{forvar259}) ?
                  reg334 : reg297)));
        end
    end
  assign wire362 = $signed($signed($unsigned((reg231[(4'h8):(1'h1)] ?
                       (^~(8'ha7)) : reg208))));
  assign wire363 = reg228;
  assign wire364 = "Fn4";
  always
    @(posedge clk) begin
      for (forvar365 = (1'h0); (forvar365 < (2'h3)); forvar365 = (forvar365 + (1'h1)))
        begin
          for (forvar366 = (1'h0); (forvar366 < (2'h2)); forvar366 = (forvar366 + (1'h1)))
            begin
              reg367 <= reg282;
              reg368 <= {$unsigned($unsigned(((-reg227) <= (reg301 ?
                      (8'ha5) : forvar314)))),
                  $unsigned({$unsigned((~^(8'ha4))), reg311})};
              reg369 = forvar280;
              reg370 = reg212[(2'h3):(2'h2)];
            end
        end
      for (forvar371 = (1'h0); (forvar371 < (2'h3)); forvar371 = (forvar371 + (1'h1)))
        begin
          reg372 <= {(7'h42)};
          for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
            begin
              reg374 = $signed($signed(("" ?
                  (~|(reg361 >> reg295)) : $signed((^reg234)))));
              reg375 <= $unsigned(reg275[(4'h9):(4'h9)]);
            end
          reg376 <= ((reg273 < (reg283[(4'hc):(4'h8)] >>> ((reg358 ?
                  (8'ha5) : (8'h9f)) ?
              $unsigned(reg329) : (reg337 ? reg316 : reg263)))) >> reg319);
          for (forvar377 = (1'h0); (forvar377 < (1'h0)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 = $unsigned((-$unsigned(((~&wire205) ?
                  $signed(reg341) : (8'hbc)))));
            end
        end
    end
  assign wire379 = forvar340;
  always
    @(posedge clk) begin
      reg380 <= (&{(((~wire239) ?
              $unsigned(reg349) : reg212[(2'h3):(1'h0)]) - forvar229)});
      if ($signed((8'ha8)))
        begin
          if (wire204[(2'h2):(1'h0)])
            begin
              reg381 = ($signed({reg331,
                  $unsigned((forvar226 ~^ reg315))}) <<< {((wire203 ?
                      "aJ4QRPucl9U09q" : forvar221) == reg272)});
            end
          else
            begin
              reg381 = (8'ha1);
              reg382 <= (!(($unsigned(wire200[(2'h2):(2'h2)]) << $unsigned({reg209})) << (~&((wire240 ?
                  reg264 : forvar371) && $signed(reg334)))));
            end
          for (forvar383 = (1'h0); (forvar383 < (1'h0)); forvar383 = (forvar383 + (1'h1)))
            begin
              reg384 <= {(reg258[(1'h0):(1'h0)] ?
                      ($signed({reg244, forvar309}) | ({(8'had)} ?
                          "CLqqL3aoEYMn" : (reg359 ?
                              forvar310 : forvar377))) : ((~&reg346[(1'h1):(1'h1)]) ?
                          forvar373 : $signed("VLfYS3UkI7giT5K9Ga"))),
                  $unsigned((8'ha9))};
              reg385 <= $signed(($signed($unsigned($signed(forvar220))) ?
                  $signed($unsigned($unsigned(reg306))) : ({{reg368, reg307},
                          (~reg342)} ?
                      (~reg315) : reg375[(4'hd):(4'hc)])));
              reg386 <= (wire362[(4'hb):(4'hb)] ?
                  forvar377 : ((($unsigned(reg316) ?
                          {reg234} : reg346) - $signed({(8'haa), reg298})) ?
                      ($signed((reg342 ^~ forvar241)) ?
                          (reg254 == reg225[(1'h1):(1'h0)]) : reg286[(5'h12):(4'he)]) : reg248));
              reg387 = (^(+$unsigned($unsigned({(8'hb4), reg306}))));
            end
          for (forvar388 = (1'h0); (forvar388 < (2'h2)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 = (~(reg278 ^ $signed($signed((wire200 ?
                  reg320 : forvar230)))));
              reg390 <= ($unsigned(((|(reg228 ? reg214 : reg295)) ?
                  (wire203[(3'h5):(1'h0)] < ((7'h42) ~^ reg231)) : $unsigned($unsigned(reg210)))) - reg386);
              reg391 <= $unsigned($unsigned((|reg387[(4'hf):(1'h0)])));
              reg392 = (^(!forvar259));
            end
          reg393 <= (reg370[(4'h8):(3'h5)] ? $signed("aW0") : (7'h44));
          reg394 <= reg353;
        end
      else
        begin
          if ({({($signed(forvar220) ?
                      reg256 : (!(8'haf)))} ^~ {reg335[(3'h4):(2'h3)],
                  (reg256 ^ $unsigned(reg337))})})
            begin
              reg381 = $signed(($signed({reg337,
                  (~&reg211)}) <<< (reg381[(2'h3):(2'h2)] > {forvar229[(2'h2):(2'h2)],
                  $unsigned(reg222)})));
              reg382 = $unsigned((reg234 && ((^~reg254) ?
                  $unsigned($unsigned(forvar351)) : reg337[(3'h4):(2'h3)])));
              reg383 <= reg271[(3'h4):(2'h2)];
              reg384 = (~$unsigned(({$unsigned(reg245), {reg344}} ?
                  (^~$unsigned(reg312)) : (reg244 >> (!(8'hb7))))));
            end
          else
            begin
              reg381 <= reg303;
              reg382 = ((~|forvar261) ^ $unsigned(((reg338 ?
                  {reg308} : (~|reg391)) <= (reg276 ?
                  reg210 : (reg215 != forvar226)))));
              reg383 = forvar310[(3'h6):(3'h6)];
            end
          reg385 = (~|($unsigned(forvar310[(3'h4):(1'h0)]) ~^ (((reg291 ?
                  reg290 : wire332) ?
              (reg387 && reg348) : $unsigned(reg245)) ^ wire364[(1'h1):(1'h1)])));
          for (forvar386 = (1'h0); (forvar386 < (2'h3)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 = forvar294[(3'h4):(1'h0)];
              reg388 <= (reg287[(5'h13):(4'hb)] >= $signed(reg246));
              reg389 = reg331;
              reg390 = (~&(8'hb7));
              reg391 = $unsigned(wire204[(3'h4):(2'h3)]);
            end
        end
      reg395 = ((8'ha7) ? wire202 : (^(reg214 << (^reg275[(3'h6):(2'h2)]))));
      reg396 <= $unsigned(forvar226);
      if ((^~$unsigned($signed($unsigned(((8'ha9) ~^ reg303))))))
        begin
          reg397 <= $unsigned(((($unsigned(wire204) ^ wire363) ^~ reg271) > (~&(&$signed(reg388)))));
        end
      else
        begin
          if ((8'hb0))
            begin
              reg397 <= forvar220;
              reg398 <= forvar377;
              reg399 <= $unsigned($unsigned((-(reg345 ^ {reg367}))));
              reg400 <= $unsigned(($signed(((reg231 << (8'ha3)) + (forvar310 ?
                      reg256 : forvar288))) ?
                  {(&(~&reg294))} : forvar347));
              reg401 = (reg246 ?
                  $unsigned((+$signed((reg258 ?
                      (8'hb3) : wire202)))) : reg376[(2'h3):(1'h0)]);
            end
          else
            begin
              reg397 = reg219;
              reg398 <= {reg254[(3'h4):(1'h0)], reg212};
              reg399 = $signed(reg250[(1'h1):(1'h0)]);
            end
          reg402 <= (~$signed(reg353[(2'h2):(1'h1)]));
          if (({wire240, (&$signed((forvar233 >>> reg345)))} ?
              $unsigned({$signed("RsXeEEDvZ0QNJo7yd"),
                  forvar322[(2'h3):(1'h0)]}) : reg393[(3'h4):(3'h4)]))
            begin
              reg403 <= (-$signed($signed({reg346[(4'hc):(4'hb)]})));
              reg404 = (-reg388);
              reg405 = {forvar383};
              reg406 <= (reg273 ?
                  ($unsigned((&reg327[(4'hf):(2'h2)])) ?
                      reg397[(2'h2):(1'h0)] : $signed(($unsigned((8'hb0)) & $unsigned(forvar340)))) : ((~^$unsigned(((8'haa) | reg385))) + forvar230[(2'h3):(2'h3)]));
            end
          else
            begin
              reg403 <= reg219[(5'h11):(2'h2)];
              reg404 = reg400[(1'h0):(1'h0)];
              reg405 <= wire200[(1'h1):(1'h1)];
              reg406 <= $unsigned(forvar269[(3'h6):(1'h0)]);
            end
          reg407 <= reg393;
        end
    end
  assign wire408 = $signed($unsigned((8'had)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module82
#( parameter param195 = {((&{{(8'h9d), (8'hbd)}}) ? ((((8'h9f) ? (8'ha8) : (8'had)) ? ((7'h41) == (7'h44)) : ((8'hb2) ? (8'ha1) : (7'h40))) ? (((8'hb8) ? (8'h9d) : (8'hbe)) << ((8'ha0) >= (7'h41))) : {((7'h44) ? (8'ha6) : (8'hba))}) : {(((8'hbe) >= (8'ha5)) + {(8'ha5)}), (((8'hb7) ? (8'h9c) : (8'hba)) > ((8'hb4) | (8'ha5)))})}
, parameter param196 = ((^~((8'haa) ? ((param195 ? param195 : param195) >> (-param195)) : (~(param195 ? param195 : (7'h44))))) >= (((8'hb3) ^~ ((param195 ? param195 : (8'haa)) & param195)) ? (^({(8'hb1)} <= (^param195))) : {(~&param195), {(param195 ? param195 : param195), (param195 >= param195)}})) )
(y, clk, wire87, wire86, wire85, wire84, wire83);
  output wire [(32'h499):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire87;
  input wire [(4'hc):(1'h0)] wire86;
  input wire [(4'hf):(1'h0)] wire85;
  input wire signed [(2'h3):(1'h0)] wire84;
  input wire [(4'hf):(1'h0)] wire83;
  wire [(3'h7):(1'h0)] wire194;
  reg [(4'hf):(1'h0)] reg193 = (1'h0);
  reg [(4'hf):(1'h0)] reg192 = (1'h0);
  reg [(4'hf):(1'h0)] reg191 = (1'h0);
  reg [(5'h15):(1'h0)] reg190 = (1'h0);
  reg [(3'h4):(1'h0)] reg189 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar188 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg187 = (1'h0);
  reg [(3'h6):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(5'h11):(1'h0)] reg182 = (1'h0);
  reg [(4'hf):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg180 = (1'h0);
  reg [(4'hb):(1'h0)] reg179 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg178 = (1'h0);
  reg [(2'h3):(1'h0)] forvar177 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg176 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg174 = (1'h0);
  reg [(4'hc):(1'h0)] reg173 = (1'h0);
  reg [(4'hc):(1'h0)] reg172 = (1'h0);
  reg [(5'h13):(1'h0)] forvar171 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar170 = (1'h0);
  reg [(4'h8):(1'h0)] reg169 = (1'h0);
  reg [(5'h15):(1'h0)] reg168 = (1'h0);
  wire [(4'he):(1'h0)] wire167;
  reg [(3'h5):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg164 = (1'h0);
  reg [(5'h11):(1'h0)] reg163 = (1'h0);
  reg [(4'he):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar160 = (1'h0);
  reg [(5'h10):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg158 = (1'h0);
  reg [(2'h2):(1'h0)] reg157 = (1'h0);
  reg [(2'h2):(1'h0)] reg156 = (1'h0);
  reg [(2'h2):(1'h0)] forvar155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg152 = (1'h0);
  reg [(3'h7):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar150 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg149 = (1'h0);
  reg [(3'h4):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg [(4'hc):(1'h0)] forvar146 = (1'h0);
  reg [(4'hc):(1'h0)] forvar145 = (1'h0);
  reg [(5'h13):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg143 = (1'h0);
  reg [(3'h5):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar139 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg138 = (1'h0);
  reg [(3'h4):(1'h0)] forvar134 = (1'h0);
  reg [(5'h15):(1'h0)] reg137 = (1'h0);
  reg [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(3'h5):(1'h0)] reg135 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg134 = (1'h0);
  wire [(5'h10):(1'h0)] wire133;
  wire signed [(5'h13):(1'h0)] wire132;
  wire signed [(5'h13):(1'h0)] wire131;
  reg [(4'hd):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg129 = (1'h0);
  reg [(3'h4):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg127 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar126 = (1'h0);
  reg [(5'h15):(1'h0)] reg125 = (1'h0);
  reg [(2'h3):(1'h0)] reg124 = (1'h0);
  reg [(3'h5):(1'h0)] reg123 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar121 = (1'h0);
  reg [(3'h5):(1'h0)] forvar120 = (1'h0);
  wire [(4'hf):(1'h0)] wire119;
  reg [(4'h8):(1'h0)] reg118 = (1'h0);
  reg [(5'h14):(1'h0)] reg117 = (1'h0);
  reg [(5'h10):(1'h0)] reg116 = (1'h0);
  reg [(5'h11):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg113 = (1'h0);
  reg [(4'he):(1'h0)] forvar112 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg111 = (1'h0);
  reg [(4'hb):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar109 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg107 = (1'h0);
  reg [(5'h13):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg105 = (1'h0);
  reg [(4'ha):(1'h0)] reg104 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar103 = (1'h0);
  reg [(4'hc):(1'h0)] reg102 = (1'h0);
  reg [(2'h3):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar100 = (1'h0);
  reg [(5'h12):(1'h0)] forvar99 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg97 = (1'h0);
  reg [(4'h8):(1'h0)] forvar96 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg95 = (1'h0);
  reg [(3'h6):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg93 = (1'h0);
  reg [(5'h14):(1'h0)] reg92 = (1'h0);
  reg [(4'ha):(1'h0)] reg91 = (1'h0);
  reg [(2'h3):(1'h0)] forvar90 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire89;
  wire [(5'h10):(1'h0)] wire88;
  assign y = {wire194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 forvar188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 forvar177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 forvar171,
                 forvar170,
                 reg169,
                 reg168,
                 wire167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 forvar160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 forvar155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 forvar150,
                 reg149,
                 reg148,
                 reg147,
                 forvar146,
                 forvar145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 forvar139,
                 reg138,
                 forvar134,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 wire133,
                 wire132,
                 wire131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 forvar126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 forvar120,
                 wire119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg110,
                 forvar109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 forvar103,
                 reg102,
                 reg101,
                 forvar100,
                 forvar99,
                 reg98,
                 reg97,
                 forvar96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 forvar90,
                 wire89,
                 wire88,
                 (1'h0)};
  assign wire88 = wire85[(3'h4):(3'h4)];
  assign wire89 = wire84;
  always
    @(posedge clk) begin
      for (forvar90 = (1'h0); (forvar90 < (2'h2)); forvar90 = (forvar90 + (1'h1)))
        begin
          if (wire86[(3'h7):(1'h0)])
            begin
              reg91 = $unsigned($signed((|{(wire85 == wire89), wire87})));
              reg92 <= $signed($unsigned((({wire84, wire86} ?
                      (~|(8'h9d)) : $signed(reg91)) ?
                  ((|(8'ha8)) ^ $unsigned(wire87)) : {$signed(wire83),
                      wire87[(4'hd):(3'h6)]})));
              reg93 <= wire85;
              reg94 <= {reg91};
              reg95 <= (!($signed((~&wire84[(2'h3):(2'h2)])) ?
                  wire83 : ((~(forvar90 & wire88)) ?
                      (~|(wire87 ? wire85 : (8'hbf))) : ("KI0" * (|wire88)))));
            end
          else
            begin
              reg91 = $signed(reg93[(2'h2):(2'h2)]);
              reg92 = reg91[(2'h2):(1'h1)];
            end
          for (forvar96 = (1'h0); (forvar96 < (2'h3)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 <= wire89;
              reg98 <= (8'h9c);
            end
        end
      for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
        begin
          for (forvar100 = (1'h0); (forvar100 < (1'h1)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 <= (((!$signed((reg97 ^~ wire83))) ?
                  forvar100[(2'h2):(1'h1)] : $signed($signed(reg91[(2'h3):(2'h2)]))) ^~ wire83);
              reg102 <= $signed(($signed($signed((reg93 | forvar90))) ^~ (((wire84 != forvar96) ?
                      {reg101, forvar99} : reg97[(3'h4):(1'h1)]) ?
                  (|(wire87 * (8'hbc))) : ((|reg98) != $signed(forvar100)))));
            end
          for (forvar103 = (1'h0); (forvar103 < (2'h3)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 <= (|$unsigned(forvar90));
              reg105 = ((forvar96 > forvar96) ?
                  (8'ha5) : $unsigned({reg91, {reg95[(1'h0):(1'h0)], wire85}}));
              reg106 <= (8'ha7);
              reg107 <= reg106;
            end
          reg108 <= wire86;
          for (forvar109 = (1'h0); (forvar109 < (1'h0)); forvar109 = (forvar109 + (1'h1)))
            begin
              reg110 = {reg95[(3'h4):(2'h3)], reg97[(1'h1):(1'h0)]};
              reg111 = "sJJd1QLAr7";
            end
          for (forvar112 = (1'h0); (forvar112 < (1'h0)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= reg107[(1'h0):(1'h0)];
              reg114 <= (^~($unsigned(((reg101 * wire84) != {wire86})) ?
                  (-(reg101[(1'h0):(1'h0)] ?
                      reg98[(4'hb):(3'h5)] : (^~(8'ha8)))) : reg93[(4'h8):(1'h0)]));
              reg115 = (+forvar100);
              reg116 = (reg101 != reg91[(1'h0):(1'h0)]);
              reg117 <= ({$signed((reg102 * (wire83 <= reg93)))} < $unsigned((8'ha4)));
            end
        end
      reg118 <= {(+((~|reg114[(2'h2):(1'h1)]) - reg117[(3'h4):(2'h3)])),
          $unsigned((^((forvar112 < (8'hac)) ? $unsigned(reg95) : reg108)))};
    end
  assign wire119 = reg102;
  always
    @(posedge clk) begin
      for (forvar120 = (1'h0); (forvar120 < (3'h4)); forvar120 = (forvar120 + (1'h1)))
        begin
          for (forvar121 = (1'h0); (forvar121 < (2'h3)); forvar121 = (forvar121 + (1'h1)))
            begin
              reg122 = reg98;
            end
          if ((~&reg97))
            begin
              reg123 <= wire83[(4'h9):(1'h1)];
              reg124 = ((-forvar99[(5'h11):(5'h10)]) >> $unsigned(({(~&forvar103)} ?
                  ((!reg95) ? (8'hbf) : $signed(wire84)) : "mEtFglEVSOY")));
            end
          else
            begin
              reg123 <= (|($unsigned(({reg94, reg92} ?
                  (wire83 ? wire83 : reg98) : (forvar96 ?
                      forvar99 : wire85))) << (~^$signed(forvar109))));
              reg124 <= (!"OVp0X2LApKu3");
              reg125 <= ((^(reg122 | (8'hbc))) == $unsigned(reg94));
            end
          for (forvar126 = (1'h0); (forvar126 < (2'h3)); forvar126 = (forvar126 + (1'h1)))
            begin
              reg127 <= (reg114[(1'h0):(1'h0)] ?
                  $signed((+((reg116 ?
                      (8'hb9) : wire87) ^~ $signed((8'hb8))))) : ((~|((wire84 ?
                      wire88 : (7'h40)) || (~reg106))) != wire89[(3'h5):(3'h4)]));
              reg128 <= (+(reg105 >>> $unsigned({(wire86 ?
                      reg107 : (8'hb2))})));
              reg129 <= (forvar126[(2'h2):(1'h0)] ?
                  ((8'hb8) && (wire86 | reg117)) : $unsigned((((+wire88) >= (reg92 ?
                          reg95 : forvar112)) ?
                      $unsigned((reg111 == (8'hba))) : reg93)));
            end
          reg130 = reg105;
        end
    end
  assign wire131 = forvar112;
  assign wire132 = ($unsigned((~^($unsigned(forvar112) ?
                           (&reg104) : ((8'hab) | forvar126)))) ?
                       {(((~|reg102) || forvar90) | (reg122[(1'h0):(1'h0)] ~^ reg107[(2'h2):(1'h1)]))} : $unsigned($signed(reg108[(1'h0):(1'h0)])));
  assign wire133 = reg123[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      if ((((^$unsigned((forvar103 ? reg111 : reg94))) + (reg130 ?
              (^(^~wire131)) : $signed({forvar121, reg129}))) ?
          reg127[(1'h1):(1'h1)] : ((-reg114) * (~^$unsigned((reg125 && wire85))))))
        begin
          reg134 <= {forvar126[(1'h0):(1'h0)]};
          if (wire84[(2'h2):(1'h0)])
            begin
              reg135 = forvar126;
              reg136 = reg128[(2'h3):(1'h1)];
            end
          else
            begin
              reg135 = $signed(reg98[(5'h12):(4'h8)]);
              reg136 = (wire131 * (reg102[(3'h7):(1'h0)] ?
                  $unsigned($signed("Qwtx2pr")) : (~(+(|reg107)))));
              reg137 = $unsigned({(reg93 & ($unsigned(forvar109) <= (reg95 >= forvar99))),
                  $unsigned(forvar112[(4'he):(1'h1)])});
            end
        end
      else
        begin
          for (forvar134 = (1'h0); (forvar134 < (1'h0)); forvar134 = (forvar134 + (1'h1)))
            begin
              reg135 <= reg94[(1'h1):(1'h1)];
              reg136 <= wire85[(4'h9):(3'h4)];
            end
        end
      reg138 <= {((($unsigned(wire131) ? wire84[(2'h2):(1'h0)] : wire119) ?
                  ({wire131} + $unsigned((8'hb4))) : {(reg115 ?
                          reg113 : forvar120)}) ?
              (~&reg137) : (&("z8Lu" && $signed(forvar109))))};
    end
  always
    @(posedge clk) begin
      for (forvar139 = (1'h0); (forvar139 < (1'h0)); forvar139 = (forvar139 + (1'h1)))
        begin
          if (reg136)
            begin
              reg140 <= reg94[(2'h3):(2'h2)];
              reg141 <= {forvar126[(1'h1):(1'h0)],
                  {$unsigned({$signed(forvar120)}),
                      (($signed(reg98) ?
                          (forvar103 <= reg97) : (reg135 ?
                              reg114 : reg107)) >> $signed((wire87 != wire87)))}};
              reg142 <= reg105[(2'h2):(1'h1)];
              reg143 <= {($signed(((~^reg104) ?
                      $unsigned(reg127) : {reg118, reg106})) <<< {{(reg93 ?
                              reg104 : reg135)},
                      (~|$signed(forvar109))})};
              reg144 <= $unsigned("RXKbhoMy");
            end
          else
            begin
              reg140 <= "9tIs1SAQX8126rr7";
              reg141 = forvar109;
              reg142 <= $signed($unsigned({wire88[(3'h5):(1'h1)],
                  (!(+reg104))}));
              reg143 <= ($unsigned($unsigned((~((8'haf) <= (8'hab))))) ?
                  reg93 : (forvar134[(2'h2):(2'h2)] ?
                      ((reg114 * reg127[(1'h1):(1'h0)]) ?
                          $signed($signed((8'ha2))) : forvar100[(4'hb):(2'h2)]) : $signed(($unsigned(wire87) ?
                          (&forvar96) : (!reg136)))));
              reg144 <= (+$signed(("kQh2zLHIcWX" ~^ ($unsigned(reg106) >>> wire132))));
            end
        end
      for (forvar145 = (1'h0); (forvar145 < (1'h0)); forvar145 = (forvar145 + (1'h1)))
        begin
          for (forvar146 = (1'h0); (forvar146 < (1'h0)); forvar146 = (forvar146 + (1'h1)))
            begin
              reg147 <= wire86[(4'h8):(1'h0)];
              reg148 <= $signed($unsigned(reg141));
              reg149 <= (|$signed(reg105));
            end
          for (forvar150 = (1'h0); (forvar150 < (3'h4)); forvar150 = (forvar150 + (1'h1)))
            begin
              reg151 = (^(~|(-(8'hbb))));
              reg152 = {reg148,
                  (wire119[(4'h8):(3'h7)] ?
                      (((reg108 ? reg92 : reg110) << (reg105 ?
                              reg147 : wire132)) ?
                          $unsigned($signed((7'h40))) : reg92[(3'h4):(1'h0)]) : (wire83 ?
                          ((forvar112 ? reg140 : reg122) ?
                              forvar103 : ((8'hbf) ?
                                  reg98 : reg108)) : forvar145[(3'h4):(1'h0)]))};
              reg153 <= reg91;
            end
          reg154 = (reg149 ?
              $signed($signed({reg115[(5'h10):(3'h5)],
                  reg92[(1'h0):(1'h0)]})) : forvar120);
          for (forvar155 = (1'h0); (forvar155 < (3'h4)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 <= {$signed(({(wire89 ? (8'hae) : (8'ha3)),
                          (^~forvar139)} ?
                      {(reg107 || wire86)} : (wire131[(3'h5):(3'h4)] ?
                          $unsigned(reg124) : (wire131 && reg129)))),
                  reg92[(4'h8):(2'h2)]};
              reg157 = $signed(($signed($signed({reg92})) > {((forvar100 ?
                          reg92 : forvar145) ?
                      (forvar90 & reg149) : $signed(reg124)),
                  $unsigned((forvar112 >>> wire132))}));
              reg158 = (^$unsigned(reg127[(1'h0):(1'h0)]));
              reg159 <= reg134;
            end
          for (forvar160 = (1'h0); (forvar160 < (3'h4)); forvar160 = (forvar160 + (1'h1)))
            begin
              reg161 = $signed((reg151 != ($signed(reg118) ?
                  ($unsigned(reg135) ?
                      (^~reg142) : (reg128 ?
                          (8'h9f) : (8'hb8))) : ($signed(reg152) != (wire89 ?
                      wire88 : reg156)))));
              reg162 = $signed((($signed({reg98,
                  wire132}) & $signed(reg92)) ^~ reg116));
              reg163 <= $unsigned($signed(($unsigned((^reg153)) - wire86[(3'h4):(1'h0)])));
              reg164 = $unsigned(reg136[(1'h0):(1'h0)]);
              reg165 = ((~^$signed((forvar121 ^ $unsigned(wire85)))) * "hR");
            end
        end
      reg166 = (8'had);
    end
  assign wire167 = ((forvar134[(2'h2):(2'h2)] | $signed(reg101[(2'h2):(1'h0)])) ?
                       reg106 : (((^~$unsigned(reg124)) ?
                           {forvar103[(3'h4):(2'h2)],
                               forvar121[(2'h2):(2'h2)]} : reg147) <<< "gL5zM93is"));
  always
    @(posedge clk) begin
      reg168 <= $unsigned(reg161[(4'hf):(1'h0)]);
      reg169 <= $unsigned({$signed(reg144[(3'h6):(3'h6)]),
          reg114[(3'h4):(1'h1)]});
      for (forvar170 = (1'h0); (forvar170 < (2'h2)); forvar170 = (forvar170 + (1'h1)))
        begin
          for (forvar171 = (1'h0); (forvar171 < (1'h0)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 <= $signed((reg97 ? (^reg137) : forvar150));
              reg173 = $unsigned((8'haf));
              reg174 = (((reg107[(1'h0):(1'h0)] == (forvar170[(3'h4):(1'h0)] ?
                      reg111 : forvar100)) ?
                  (reg159 ^~ $signed($unsigned((8'hba)))) : ($unsigned((reg105 ~^ reg114)) < ((reg142 ?
                      reg153 : reg95) | "lphJ31l7"))) + (reg148[(3'h4):(1'h0)] ?
                  wire131[(4'hb):(4'ha)] : wire131));
              reg175 <= (|(~&(!wire86)));
              reg176 = reg152[(4'he):(4'hc)];
            end
          for (forvar177 = (1'h0); (forvar177 < (2'h3)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 = $signed(reg104[(3'h7):(3'h7)]);
              reg179 <= (&(~^((reg111[(4'h8):(3'h6)] ?
                      forvar160[(5'h15):(3'h7)] : (^wire87)) ?
                  $unsigned((+(8'hae))) : (~$unsigned((8'h9d))))));
            end
          reg180 = wire131[(5'h11):(5'h10)];
          reg181 = $signed(((reg161[(1'h0):(1'h0)] ^ ((^~forvar155) ?
              forvar126[(4'h9):(3'h6)] : $unsigned(reg102))) >>> wire167));
          if ($signed((!(!($signed(reg136) <= reg134)))))
            begin
              reg182 <= reg153;
              reg183 <= $unsigned($unsigned(((&((7'h43) ?
                  wire89 : reg102)) <= (forvar139 ?
                  (reg130 ? forvar170 : forvar134) : (reg110 + reg153)))));
              reg184 <= $signed($unsigned(($signed({wire85, reg142}) ?
                  ($unsigned(forvar103) && $signed(reg122)) : reg147)));
              reg185 <= reg97;
              reg186 <= reg107[(3'h7):(2'h2)];
            end
          else
            begin
              reg182 <= ((~^forvar150[(3'h5):(3'h5)]) ?
                  reg159 : ((|wire89[(2'h3):(2'h3)]) ?
                      $signed((^~$signed(wire89))) : (~&"ZOl4NEMRZNlIz")));
              reg183 = (reg101 ?
                  $unsigned(reg108) : $unsigned($signed($signed($unsigned((8'ha2))))));
              reg184 <= wire132;
              reg185 = $unsigned($unsigned(($unsigned(reg161[(3'h4):(3'h4)]) ?
                  "5wrvG" : $unsigned($signed(reg104)))));
              reg186 <= forvar109;
            end
        end
      reg187 <= forvar109[(3'h4):(2'h2)];
      for (forvar188 = (1'h0); (forvar188 < (3'h4)); forvar188 = (forvar188 + (1'h1)))
        begin
          if (reg142)
            begin
              reg189 <= ($unsigned($signed(forvar120)) << ((~(reg186 != $unsigned(reg157))) ?
                  reg140 : ($unsigned($unsigned(forvar126)) ~^ (reg128 ?
                      reg172 : {wire86, (8'hab)}))));
              reg190 = ((((8'ha4) ~^ reg173) ?
                      (($signed((8'hbf)) | $signed(reg143)) ?
                          {$signed(reg185),
                              (wire133 ?
                                  reg187 : reg125)} : ($unsigned(reg129) ~^ {(7'h40),
                              wire86})) : (({reg113, reg116} ?
                              $unsigned(forvar139) : $signed(reg174)) ?
                          $unsigned(reg178[(2'h2):(2'h2)]) : ({forvar155} << reg149[(1'h1):(1'h0)]))) ?
                  $unsigned((!reg137[(4'hc):(3'h6)])) : reg163[(4'hf):(4'hc)]);
            end
          else
            begin
              reg189 = (|(&(|(!(reg182 ? reg122 : reg102)))));
              reg190 = reg181[(2'h3):(1'h1)];
              reg191 <= $signed({$unsigned(((8'hb5) << $signed(forvar171)))});
              reg192 = (8'ha6);
              reg193 <= $signed(wire132);
            end
        end
    end
  assign wire194 = $signed("rPe5R3O9rdG9N1");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module29
#( parameter param55 = ({(7'h41)} ? {(~|(~&{(7'h40)})), ((((8'hbc) ? (8'hb0) : (8'ha3)) ? (+(8'hbb)) : ((8'hac) < (8'hbb))) ? (8'hb1) : (&(8'hbd)))} : {((8'had) && (((8'hb5) ? (8'h9f) : (8'ha3)) ? (&(8'hb8)) : ((8'hb4) || (8'hb2)))), ((8'haf) ? {{(7'h43), (8'hbb)}} : ((+(7'h41)) || (~|(8'hb4))))})
, parameter param56 = (~|((8'ha6) <= (8'hb2))) )
(y, clk, wire33, wire32, wire31, wire30);
  output wire [(32'hc5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire33;
  input wire signed [(3'h6):(1'h0)] wire32;
  input wire signed [(4'hf):(1'h0)] wire31;
  input wire signed [(5'h10):(1'h0)] wire30;
  wire [(2'h3):(1'h0)] wire54;
  wire signed [(5'h13):(1'h0)] wire53;
  wire signed [(3'h7):(1'h0)] wire52;
  wire [(4'hb):(1'h0)] wire51;
  wire [(3'h6):(1'h0)] wire50;
  wire [(4'h8):(1'h0)] wire49;
  wire signed [(4'hd):(1'h0)] wire48;
  wire signed [(2'h3):(1'h0)] wire47;
  wire [(4'he):(1'h0)] wire46;
  wire [(3'h6):(1'h0)] wire45;
  wire signed [(4'h8):(1'h0)] wire44;
  wire signed [(4'h8):(1'h0)] wire43;
  reg [(3'h7):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg41 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg40 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar38 = (1'h0);
  reg [(5'h10):(1'h0)] forvar37 = (1'h0);
  wire [(2'h3):(1'h0)] wire36;
  wire signed [(3'h6):(1'h0)] wire35;
  wire [(4'hc):(1'h0)] wire34;
  assign y = {wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 wire48,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 forvar38,
                 forvar37,
                 wire36,
                 wire35,
                 wire34,
                 (1'h0)};
  assign wire34 = wire30;
  assign wire35 = (^~(wire33[(5'h12):(4'h8)] ^~ (~&{wire32, (-wire30)})));
  assign wire36 = wire31[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar37 = (1'h0); (forvar37 < (1'h0)); forvar37 = (forvar37 + (1'h1)))
        begin
          for (forvar38 = (1'h0); (forvar38 < (2'h2)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 = wire35;
              reg40 <= ($signed(forvar37[(4'h8):(3'h6)]) ?
                  forvar37[(3'h4):(1'h1)] : $signed($unsigned($unsigned(wire36[(1'h0):(1'h0)]))));
              reg41 = $unsigned(($signed((-(wire32 ? wire32 : reg40))) ?
                  ($unsigned($signed(reg39)) <= ({(8'ha4)} ?
                      $unsigned(forvar38) : (wire36 ?
                          forvar37 : (7'h41)))) : {wire32[(3'h4):(1'h0)]}));
            end
          reg42 <= ($signed($signed({reg40[(4'h8):(2'h3)],
                  $signed(forvar37)})) ?
              forvar37[(4'hb):(3'h4)] : $unsigned($signed($signed((wire34 ?
                  (8'h9e) : wire35)))));
        end
    end
  assign wire43 = (8'hb7);
  assign wire44 = (forvar37[(2'h3):(1'h1)] >>> (forvar38[(4'hf):(4'ha)] ?
                      $signed(forvar38[(2'h3):(2'h3)]) : wire30));
  assign wire45 = $signed($unsigned(($unsigned((!wire35)) << ($signed(reg39) > ((8'hae) ?
                      wire33 : (8'ha0))))));
  assign wire46 = "";
  assign wire47 = (|wire34);
  assign wire48 = reg42;
  assign wire49 = forvar37;
  assign wire50 = ((8'hbb) ?
                      wire44[(1'h0):(1'h0)] : {{wire47, reg42[(3'h5):(2'h3)]}});
  assign wire51 = $signed((~^wire49));
  assign wire52 = {reg42[(2'h3):(2'h3)]};
  assign wire53 = wire35;
  assign wire54 = (~|reg41);
endmodule
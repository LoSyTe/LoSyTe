(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param978 = {(~|((8'hbd) ^ (((8'hb0) ? (8'hb3) : (8'hb0)) ? ((7'h4e) >> (8'hb1)) : ((8'hb8) ? (7'h4b) : (8'hb3)))))}, 
parameter param979 = param978)
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h989):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire0;
  input wire [(2'h3):(1'h0)] wire1;
  input wire [(4'h9):(1'h0)] wire2;
  input wire [(2'h3):(1'h0)] wire3;
  input wire [(5'h13):(1'h0)] wire4;
  wire signed [(4'h8):(1'h0)] wire36;
  wire signed [(5'h16):(1'h0)] wire86;
  wire [(4'hb):(1'h0)] wire133;
  wire signed [(5'h1a):(1'h0)] wire938;
  reg signed [(5'h17):(1'h0)] reg977 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg976 = (1'h0);
  reg [(3'h5):(1'h0)] reg975 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg974 = (1'h0);
  reg [(5'h15):(1'h0)] reg973 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg972 = (1'h0);
  reg [(3'h5):(1'h0)] reg971 = (1'h0);
  reg [(5'h18):(1'h0)] reg970 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg969 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg968 = (1'h0);
  reg [(5'h19):(1'h0)] reg967 = (1'h0);
  reg [(5'h19):(1'h0)] reg966 = (1'h0);
  reg [(2'h3):(1'h0)] reg965 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg964 = (1'h0);
  reg [(4'hb):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg962 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg960 = (1'h0);
  reg [(5'h18):(1'h0)] reg959 = (1'h0);
  reg [(3'h5):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg957 = (1'h0);
  reg [(5'h14):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg955 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg954 = (1'h0);
  reg [(2'h3):(1'h0)] reg953 = (1'h0);
  reg [(5'h10):(1'h0)] reg952 = (1'h0);
  reg [(4'hb):(1'h0)] reg951 = (1'h0);
  reg [(3'h6):(1'h0)] reg950 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg949 = (1'h0);
  reg [(4'he):(1'h0)] reg948 = (1'h0);
  reg signed [(4'he):(1'h0)] reg947 = (1'h0);
  reg [(4'ha):(1'h0)] reg946 = (1'h0);
  reg [(5'h19):(1'h0)] reg945 = (1'h0);
  reg [(4'ha):(1'h0)] reg944 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg942 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg941 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg940 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5 = (1'h0);
  reg [(4'hf):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg7 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg8 = (1'h0);
  reg [(5'h14):(1'h0)] reg9 = (1'h0);
  reg [(4'hf):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg11 = (1'h0);
  reg [(3'h6):(1'h0)] reg12 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg15 = (1'h0);
  reg [(4'ha):(1'h0)] reg16 = (1'h0);
  reg [(5'h18):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg18 = (1'h0);
  reg [(4'hc):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg20 = (1'h0);
  reg [(5'h11):(1'h0)] reg21 = (1'h0);
  reg [(4'h9):(1'h0)] reg22 = (1'h0);
  reg [(4'h8):(1'h0)] reg23 = (1'h0);
  reg [(5'h19):(1'h0)] reg24 = (1'h0);
  reg [(4'hf):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg26 = (1'h0);
  reg [(4'hf):(1'h0)] reg27 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg28 = (1'h0);
  reg [(4'hf):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg31 = (1'h0);
  reg [(5'h15):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg34 = (1'h0);
  reg [(4'hb):(1'h0)] reg35 = (1'h0);
  reg [(2'h2):(1'h0)] reg37 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg39 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg41 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg42 = (1'h0);
  reg [(5'h17):(1'h0)] reg43 = (1'h0);
  reg [(4'hb):(1'h0)] reg44 = (1'h0);
  reg [(3'h5):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg48 = (1'h0);
  reg [(5'h16):(1'h0)] reg49 = (1'h0);
  reg [(5'h14):(1'h0)] reg50 = (1'h0);
  reg [(5'h12):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg52 = (1'h0);
  reg [(4'hf):(1'h0)] reg53 = (1'h0);
  reg [(5'h12):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg57 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg60 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg61 = (1'h0);
  reg [(5'h19):(1'h0)] reg62 = (1'h0);
  reg [(4'h8):(1'h0)] reg63 = (1'h0);
  reg [(4'hc):(1'h0)] reg64 = (1'h0);
  reg [(4'h9):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg67 = (1'h0);
  reg [(4'hb):(1'h0)] reg68 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg69 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg72 = (1'h0);
  reg [(5'h10):(1'h0)] reg73 = (1'h0);
  reg [(4'he):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg75 = (1'h0);
  reg [(5'h13):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg78 = (1'h0);
  reg [(4'hd):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(2'h2):(1'h0)] reg83 = (1'h0);
  reg [(4'h8):(1'h0)] reg84 = (1'h0);
  reg [(5'h18):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(3'h5):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg94 = (1'h0);
  reg [(3'h7):(1'h0)] reg95 = (1'h0);
  reg [(3'h5):(1'h0)] reg96 = (1'h0);
  reg [(5'h15):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg98 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg99 = (1'h0);
  reg [(5'h19):(1'h0)] reg100 = (1'h0);
  reg [(4'hb):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg105 = (1'h0);
  reg [(5'h10):(1'h0)] reg106 = (1'h0);
  reg [(4'ha):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg108 = (1'h0);
  reg [(5'h18):(1'h0)] reg109 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg110 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg112 = (1'h0);
  reg [(4'hb):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg114 = (1'h0);
  reg [(5'h13):(1'h0)] reg115 = (1'h0);
  reg [(4'h8):(1'h0)] reg116 = (1'h0);
  reg [(3'h7):(1'h0)] reg117 = (1'h0);
  reg [(5'h15):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg119 = (1'h0);
  reg [(4'hc):(1'h0)] reg120 = (1'h0);
  reg [(5'h11):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg122 = (1'h0);
  reg [(5'h14):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg124 = (1'h0);
  reg [(4'hf):(1'h0)] reg125 = (1'h0);
  reg [(5'h12):(1'h0)] reg126 = (1'h0);
  reg [(3'h7):(1'h0)] reg127 = (1'h0);
  reg signed [(4'he):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg130 = (1'h0);
  reg [(5'h1a):(1'h0)] reg131 = (1'h0);
  reg [(5'h19):(1'h0)] reg132 = (1'h0);
  assign y = {wire36,
                 wire86,
                 wire133,
                 wire938,
                 reg977,
                 reg976,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 reg956,
                 reg955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 reg945,
                 reg944,
                 reg943,
                 reg942,
                 reg941,
                 reg940,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 reg60,
                 reg61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 reg78,
                 reg79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 reg129,
                 reg130,
                 reg131,
                 reg132,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire3[(1'h1):(1'h1)])
        begin
          if ((((wire0 <<< wire2[(1'h0):(1'h0)]) ?
              ($signed({wire0}) ?
                  (~wire0[(1'h1):(1'h1)]) : (^~((7'h49) ?
                      (7'h41) : wire2))) : (wire2[(2'h2):(1'h0)] == (wire1[(1'h0):(1'h0)] > wire1))) > (wire4[(2'h2):(1'h0)] ?
              (($unsigned(wire4) ? (^wire3) : (&wire4)) != (wire2 ?
                  $signed(wire3) : wire3[(2'h2):(2'h2)])) : (7'h44))))
            begin
              reg5 <= ($unsigned((((wire1 ?
                  wire1 : wire0) >>> (wire2 * wire4)) || wire1)) + (8'hb9));
              reg6 <= wire4;
              reg7 <= reg5[(1'h1):(1'h1)];
            end
          else
            begin
              reg5 <= ((reg7[(5'h16):(5'h14)] ?
                  ($unsigned($unsigned(wire0)) ^ $signed($unsigned(wire2))) : $signed(wire4[(3'h5):(1'h0)])) < ((!($unsigned(wire4) ?
                  $unsigned(wire1) : reg7[(4'he):(2'h3)])) & (wire3 ?
                  {wire1[(1'h1):(1'h1)], $signed(wire4)} : {(!wire1),
                      $unsigned(wire1)})));
              reg6 <= {(~^$unsigned(($signed(wire3) < $signed(wire3)))),
                  $unsigned($unsigned($signed($signed(reg7))))};
              reg7 <= wire3[(1'h1):(1'h1)];
              reg8 <= wire0[(3'h4):(2'h3)];
              reg9 <= $unsigned((({wire4} ?
                      ($signed(reg7) * reg7[(5'h10):(3'h4)]) : (reg6[(2'h3):(2'h2)] + $unsigned((8'ha8)))) ?
                  wire2 : $signed(($signed(wire1) ?
                      reg6 : wire1[(2'h3):(2'h2)]))));
              reg10 <= ((8'ha0) ^~ (&(^~((^reg9) ? $signed(wire2) : (^reg6)))));
            end
          reg11 <= ((($signed(wire0) ?
                  (reg10[(3'h7):(3'h5)] >> wire3[(2'h2):(1'h1)]) : reg7[(3'h6):(1'h1)]) ?
              (-reg6) : $unsigned(reg8[(3'h4):(2'h2)])) + ($unsigned((^$unsigned(wire4))) >= (((~reg6) <<< $unsigned((7'h4c))) >> reg9)));
          reg12 <= reg7[(5'h17):(5'h16)];
          if ($signed((($signed((reg10 ? wire4 : wire1)) ?
                  (^$signed(wire1)) : ((reg12 != reg9) < reg8)) ?
              (7'h40) : wire0[(3'h4):(2'h2)])))
            begin
              reg13 <= (reg9 ?
                  (~$signed(reg11[(3'h5):(2'h3)])) : ($signed($unsigned(wire0[(1'h0):(1'h0)])) < $unsigned(reg8[(3'h5):(3'h4)])));
              reg14 <= wire4;
            end
          else
            begin
              reg13 <= wire0;
              reg14 <= $unsigned($signed(((~reg13[(2'h2):(1'h0)]) ?
                  ((^wire0) ? (reg7 <<< wire4) : {reg6, wire3}) : wire0)));
              reg15 <= ({(~|{(8'haa)}),
                  $unsigned((~wire2[(3'h7):(1'h0)]))} != {({(reg14 != wire1)} > $unsigned((wire3 && reg7))),
                  (~^(-reg13))});
            end
          reg16 <= ($unsigned((!$signed((^~(8'hb0))))) << ((($unsigned(wire4) * (reg5 ^ reg11)) * {$unsigned(reg6)}) || ({(reg15 ?
                  wire0 : (8'ha2)),
              (wire1 >>> reg11)} ^ (reg6[(1'h1):(1'h0)] ~^ $signed((8'ha9))))));
        end
      else
        begin
          reg5 <= $signed($unsigned((~{$unsigned(reg14)})));
          reg6 <= (7'h41);
        end
      if (reg12[(2'h3):(1'h0)])
        begin
          reg17 <= (!reg13[(3'h5):(1'h0)]);
          if ($unsigned($unsigned(wire3)))
            begin
              reg18 <= ((~(^~$signed(reg8[(1'h0):(1'h0)]))) ?
                  reg13 : ($signed({(7'h48)}) << (($unsigned(reg10) ?
                          $signed(reg14) : reg5) ?
                      $signed(reg9[(5'h14):(4'h9)]) : (~^{(8'ha9)}))));
              reg19 <= wire1[(1'h1):(1'h0)];
              reg20 <= (~&reg12);
            end
          else
            begin
              reg18 <= ((^~(-wire0)) ?
                  ({$unsigned((|wire1)), $signed((8'ha6))} ?
                      wire4[(5'h13):(4'hb)] : ($unsigned($signed(reg9)) << $signed((^~wire2)))) : (|$unsigned(wire2)));
              reg19 <= $signed(reg11);
              reg20 <= reg8[(3'h7):(3'h4)];
              reg21 <= ((8'ha5) ?
                  $signed((((reg20 ? reg19 : (8'hbf)) ?
                      $unsigned(reg15) : {reg19}) != reg8[(4'h8):(1'h1)])) : ((((-wire4) ?
                          {reg7} : (reg8 ^~ reg16)) ?
                      {wire0[(3'h4):(2'h2)]} : {reg5}) || reg9));
            end
          if (reg6)
            begin
              reg22 <= $signed(((~^$unsigned($signed((7'h4d)))) ?
                  {((~reg20) && wire2[(4'h8):(1'h1)]),
                      $signed(reg10)} : wire4));
              reg23 <= reg7;
              reg24 <= wire1;
            end
          else
            begin
              reg22 <= (^(-({(reg20 || (8'hb4)),
                  $signed(reg18)} || reg13[(4'h9):(3'h6)])));
              reg23 <= {wire2, $signed(reg21[(4'hd):(1'h1)])};
              reg24 <= (reg21[(1'h1):(1'h1)] ?
                  (~^$signed($signed($signed(wire2)))) : (^~{reg12,
                      $unsigned((+(8'h9f)))}));
              reg25 <= $signed(($unsigned(reg5[(2'h2):(1'h1)]) & reg18));
              reg26 <= (+reg11);
              reg27 <= $unsigned((reg19[(4'h9):(2'h2)] ?
                  $unsigned($unsigned($signed(wire4))) : $signed($signed(((8'ha1) ?
                      reg26 : reg12)))));
            end
          if ($unsigned((((wire4[(4'hf):(1'h0)] || (+reg27)) <= {$signed(reg19),
              (~|reg12)}) <<< reg9[(2'h3):(1'h0)])))
            begin
              reg28 <= reg17;
              reg29 <= {(8'ha9)};
              reg30 <= reg27;
            end
          else
            begin
              reg28 <= (reg11[(3'h5):(3'h5)] ?
                  $signed($unsigned((+$unsigned(wire3)))) : wire1);
              reg29 <= wire0[(1'h1):(1'h0)];
              reg30 <= (+$signed($unsigned(($signed(reg10) <= reg9[(5'h14):(3'h5)]))));
              reg31 <= reg9;
              reg32 <= (|$unsigned({$signed(((8'hbc) << reg22)),
                  (~(reg19 ? wire1 : wire0))}));
              reg33 <= reg6;
            end
          reg34 <= $unsigned(reg27[(2'h2):(1'h1)]);
          reg35 <= (($signed((reg5 ^~ {reg34, reg13})) ? (~&wire3) : wire0) ?
              reg8 : reg11[(3'h4):(1'h1)]);
        end
      else
        begin
          if (((wire0 ?
              reg35[(3'h5):(3'h5)] : ($unsigned((reg22 ? reg28 : (7'h40))) ?
                  ({reg25} ? (~reg19) : $signed(reg23)) : (reg28 ?
                      (8'hac) : wire3[(1'h1):(1'h0)]))) > (8'hb7)))
            begin
              reg17 <= (^~reg33[(3'h4):(1'h1)]);
              reg18 <= wire0;
            end
          else
            begin
              reg17 <= wire0[(2'h3):(1'h0)];
            end
          reg19 <= ((reg35 << ((8'ha2) + $unsigned($signed(wire2)))) ^~ $unsigned(reg27[(4'hc):(4'h8)]));
          reg20 <= {((&(reg25 ?
                  $signed(reg14) : reg16)) <<< {reg14[(4'h8):(4'h8)]})};
          reg21 <= $signed((reg11 ?
              (~^$unsigned(reg7)) : $signed((-$signed((8'hab))))));
          if (((reg33[(2'h3):(1'h1)] ?
              (+(reg31 == wire2)) : ($signed((+reg35)) ?
                  $signed(((8'hbf) && reg28)) : (~reg24[(5'h12):(4'hf)]))) - reg16[(1'h1):(1'h0)]))
            begin
              reg22 <= wire4[(3'h6):(1'h0)];
              reg23 <= $signed((reg24[(5'h12):(4'hc)] ?
                  ((reg17 ^ $signed(reg23)) + {(reg13 >= reg10)}) : wire0[(2'h3):(1'h0)]));
              reg24 <= reg25[(3'h7):(3'h7)];
              reg25 <= $unsigned(wire2[(3'h4):(2'h2)]);
              reg26 <= ((reg21 >>> {(|$unsigned(reg6)),
                  (~&((8'h9e) >>> reg14))}) != {reg29});
            end
          else
            begin
              reg22 <= wire3;
              reg23 <= ({reg7[(3'h6):(3'h4)],
                      $signed(((reg21 << reg29) ~^ (reg27 && reg11)))} ?
                  reg30 : (+(((|reg14) ? $signed(reg13) : reg9) ?
                      (!{reg13}) : (reg5[(1'h0):(1'h0)] ^ wire3))));
            end
          reg27 <= {(~|reg14)};
        end
    end
  assign wire36 = $unsigned(reg17[(4'he):(2'h3)]);
  always
    @(posedge clk) begin
      reg37 <= $signed({(reg20 ?
              (~|wire1[(2'h2):(1'h1)]) : $unsigned((reg20 ? wire2 : reg21)))});
      if ($signed(reg21))
        begin
          reg38 <= (!$unsigned(wire4));
          if (($signed(wire36[(1'h0):(1'h0)]) - {({reg21,
                      reg23[(3'h7):(3'h5)]} ?
                  ($signed((8'hbd)) & reg17) : {reg5, reg8[(1'h1):(1'h0)]}),
              $signed({{reg23, wire3}})}))
            begin
              reg39 <= reg11;
              reg40 <= reg7;
              reg41 <= reg34[(1'h0):(1'h0)];
              reg42 <= reg33[(4'hd):(4'hd)];
              reg43 <= ($unsigned(((|reg12) <<< (reg18 < $unsigned(wire4)))) <<< (8'h9f));
            end
          else
            begin
              reg39 <= reg39[(3'h4):(2'h3)];
            end
          reg44 <= $signed((~$signed(((^~reg20) && {reg19}))));
          if ($signed(reg41[(5'h11):(4'hb)]))
            begin
              reg45 <= ($signed(reg25[(1'h1):(1'h1)]) ? reg12 : wire0);
              reg46 <= reg32[(2'h3):(2'h3)];
              reg47 <= reg8[(4'h8):(3'h6)];
              reg48 <= $signed(wire2);
              reg49 <= {(~^($signed(reg9[(4'he):(1'h1)]) | $unsigned(reg8[(3'h5):(1'h0)]))),
                  (-(~&(reg48[(5'h13):(3'h7)] & (wire3 ? wire2 : reg47))))};
              reg50 <= $signed(reg41[(4'hb):(1'h1)]);
            end
          else
            begin
              reg45 <= $unsigned($signed(reg14));
              reg46 <= reg42;
              reg47 <= reg48[(4'hc):(4'hb)];
              reg48 <= reg26[(4'hc):(3'h7)];
            end
        end
      else
        begin
          reg38 <= $unsigned($signed((wire1[(2'h2):(2'h2)] + (reg32[(1'h0):(1'h0)] * (reg16 ?
              wire0 : reg14)))));
          if (reg31)
            begin
              reg39 <= reg19[(3'h7):(3'h7)];
              reg40 <= ($unsigned(($signed((~&reg27)) > (^(reg19 ?
                  (7'h46) : reg23)))) && $signed((reg48[(3'h6):(2'h3)] ?
                  {(wire4 ? reg40 : reg44), wire36} : ({reg44, (7'h46)} ?
                      (reg6 | (8'hb3)) : reg49))));
              reg41 <= {reg35};
              reg42 <= reg48;
            end
          else
            begin
              reg39 <= reg16[(4'ha):(1'h0)];
              reg40 <= reg38;
              reg41 <= (^$unsigned($signed(wire4)));
            end
          if ((~^$unsigned($unsigned(((reg10 + reg43) ?
              (reg9 < reg50) : {reg44, (7'h4d)})))))
            begin
              reg43 <= (^$signed((~&(|(reg29 ^~ reg16)))));
              reg44 <= (reg26[(3'h4):(2'h2)] ?
                  reg42 : (-(wire36 < (reg32[(4'ha):(1'h1)] ?
                      reg20 : (7'h47)))));
              reg45 <= {(|reg5[(1'h0):(1'h0)]),
                  (reg26 != (+(~&(reg12 ? wire36 : reg30))))};
              reg46 <= reg21[(2'h3):(1'h0)];
              reg47 <= {((reg19 ^ reg9[(3'h7):(3'h5)]) - reg26[(3'h5):(2'h2)])};
            end
          else
            begin
              reg43 <= reg27[(1'h1):(1'h1)];
              reg44 <= $unsigned($unsigned($unsigned(($signed(reg18) ?
                  reg23 : reg25[(4'h9):(2'h2)]))));
              reg45 <= $unsigned(wire2[(3'h4):(1'h0)]);
              reg46 <= $signed((($signed((reg11 ? reg47 : reg50)) <<< (wire2 ?
                      wire36 : (!(7'h42)))) ?
                  (+((+(8'hac)) ^~ (&wire2))) : $unsigned((-$signed(wire1)))));
              reg47 <= $signed(reg31);
              reg48 <= (!($unsigned((-$signed(reg17))) ?
                  reg38[(4'h8):(3'h5)] : wire36));
            end
          reg49 <= reg34[(4'ha):(1'h1)];
          if (($signed(reg11[(2'h3):(2'h3)]) <<< ($signed(((|reg25) < (reg27 >>> wire3))) ^ ((wire0[(3'h4):(1'h0)] ?
              $unsigned(reg47) : (reg15 ?
                  wire1 : reg14)) >= $unsigned(reg39[(3'h4):(1'h0)])))))
            begin
              reg50 <= wire4;
            end
          else
            begin
              reg50 <= reg35;
              reg51 <= $signed(reg7);
              reg52 <= {$signed(wire1),
                  $unsigned((~^($signed(reg28) ?
                      $signed(reg7) : (reg33 ? reg37 : wire0))))};
              reg53 <= wire1[(2'h2):(1'h0)];
              reg54 <= {reg39, ($unsigned(reg24) || $unsigned(reg47))};
              reg55 <= reg53[(4'hb):(3'h7)];
            end
          if (((~|$unsigned($unsigned($signed(reg50)))) ^~ $unsigned(((reg32[(5'h11):(4'hf)] ?
                  (-reg43) : {(8'h9d)}) ?
              $unsigned($signed(reg12)) : $unsigned((-reg51))))))
            begin
              reg56 <= (reg42[(1'h1):(1'h1)] <<< reg16[(4'ha):(1'h1)]);
              reg57 <= reg43[(4'h8):(3'h5)];
              reg58 <= reg30;
            end
          else
            begin
              reg56 <= reg11[(1'h0):(1'h0)];
              reg57 <= (~|(-$signed(($unsigned(reg19) - ((8'ha1) ?
                  reg48 : wire2)))));
            end
        end
      reg59 <= ($signed((8'hb8)) ?
          $signed((+((reg20 ?
              (8'hb7) : wire0) << reg8[(3'h5):(1'h1)]))) : $signed((8'ha8)));
      if (reg52)
        begin
          if ($unsigned({((|$signed(wire0)) ?
                  ((~|(7'h4a)) ?
                      reg21[(1'h0):(1'h0)] : $unsigned(reg31)) : ($unsigned(reg18) + (reg43 ?
                      (7'h47) : reg46)))}))
            begin
              reg60 <= (reg33 ?
                  $unsigned((($signed((7'h46)) & {reg41, (7'h4d)}) ?
                      ((~^wire36) < $signed(reg30)) : reg18[(4'ha):(3'h6)])) : {(8'hb4)});
              reg61 <= (~^(reg59[(4'h8):(2'h3)] ?
                  reg54 : ((^$unsigned(reg19)) >> $signed((reg11 ?
                      reg33 : reg44)))));
              reg62 <= reg5;
            end
          else
            begin
              reg60 <= reg30;
              reg61 <= ($signed((~$signed(reg21[(3'h4):(2'h2)]))) >= $unsigned((((reg37 ~^ reg40) ?
                      reg48[(1'h0):(1'h0)] : (reg18 ? reg30 : reg13)) ?
                  ({reg48} ? $signed((8'h9d)) : $signed(reg38)) : (7'h41))));
            end
          if (($unsigned($signed(((wire36 >= reg12) ?
                  reg28[(2'h3):(1'h0)] : (reg62 ? reg37 : (8'ha2))))) ?
              (-$unsigned((!reg23))) : (7'h48)))
            begin
              reg63 <= $signed({(^~($signed(reg13) ^ reg6)),
                  ($signed((reg50 < reg39)) ?
                      ((reg56 == reg24) << (7'h4c)) : (~reg22))});
            end
          else
            begin
              reg63 <= reg25[(4'hb):(4'hb)];
              reg64 <= $signed((~|($signed(reg56) ?
                  $unsigned(reg58[(4'h8):(1'h1)]) : reg56)));
            end
          reg65 <= ((wire0[(1'h0):(1'h0)] <= ($signed(reg62[(1'h0):(1'h0)]) ^ reg30[(4'hb):(3'h4)])) ?
              (~^$signed(reg26)) : (!(reg25[(3'h5):(3'h4)] ?
                  $unsigned($unsigned(reg27)) : ({wire2, reg48} ?
                      $signed((8'hb9)) : (~wire4)))));
          if ($unsigned($unsigned(reg9[(2'h2):(1'h0)])))
            begin
              reg66 <= ((+reg35) >> (~^$signed((~&reg61))));
              reg67 <= (~^((+wire1[(2'h3):(2'h3)]) ?
                  $signed(((reg28 ? reg60 : reg17) ?
                      (reg23 ? (8'hb7) : (8'h9e)) : {reg48,
                          wire0})) : (reg38[(1'h1):(1'h0)] ?
                      reg7 : {$signed(reg21)})));
              reg68 <= ($unsigned($signed($unsigned({wire36}))) ?
                  (|$signed($unsigned((reg23 ?
                      reg8 : reg58)))) : $signed($signed(wire0)));
              reg69 <= {$unsigned((+((reg28 <= reg16) | reg57)))};
              reg70 <= $signed((reg34 ?
                  {reg62[(1'h1):(1'h1)],
                      (reg34 < reg42[(1'h1):(1'h1)])} : (^~($signed(reg38) ?
                      reg26[(3'h6):(3'h4)] : wire4))));
              reg71 <= ($unsigned((+$unsigned(reg30[(3'h7):(3'h6)]))) ?
                  {{$unsigned((^~reg42)),
                          $unsigned(((7'h4b) ?
                              reg47 : wire0))}} : (+$unsigned(($signed(reg22) <= wire4[(5'h10):(2'h2)]))));
            end
          else
            begin
              reg66 <= $unsigned((~^$signed(((reg41 ?
                  reg63 : reg21) | reg59))));
              reg67 <= (((((reg39 && reg10) == reg19) ?
                      reg29 : $signed(reg12)) > $signed((-$unsigned(reg5)))) ?
                  (~|$signed(($signed(reg68) | $signed(reg45)))) : ($signed($unsigned($unsigned(reg29))) >= reg58[(3'h5):(2'h3)]));
              reg68 <= $signed((((^~(reg41 <= reg33)) ?
                  $signed($signed(reg14)) : (((8'ha2) ? reg11 : reg59) ?
                      {reg34} : $unsigned(reg30))) ^~ reg22));
              reg69 <= $signed((({(~|reg68)} ?
                  reg59 : $unsigned($signed(reg64))) <<< $unsigned(($unsigned(wire3) << (reg27 ?
                  reg42 : reg66)))));
            end
        end
      else
        begin
          if ({{wire4, reg45[(1'h0):(1'h0)]},
              ((8'ha5) || {reg13[(4'hb):(2'h2)]})})
            begin
              reg60 <= (($signed($unsigned((reg39 + reg23))) ?
                      $unsigned(reg41) : $signed($unsigned($signed(reg47)))) ?
                  (({reg46, $unsigned(reg54)} ^~ reg40[(4'hb):(3'h7)]) ?
                      ($unsigned($unsigned(reg29)) ?
                          ((^~reg50) && $signed((8'ha0))) : reg21[(4'he):(4'h8)]) : reg68) : ({$unsigned($signed(reg31))} <= (!$signed(reg52[(5'h14):(4'hf)]))));
            end
          else
            begin
              reg60 <= ($unsigned($unsigned(((&(8'hb5)) ?
                  reg61 : {reg61, reg55}))) ^~ (reg61 ?
                  (^~(^~(^~reg60))) : ((+(reg23 == reg30)) ?
                      reg54[(4'h8):(1'h1)] : reg58)));
            end
        end
      if ($signed(reg53[(4'he):(3'h7)]))
        begin
          if (reg5)
            begin
              reg72 <= (~reg71);
            end
          else
            begin
              reg72 <= $unsigned(((7'h43) > {$signed($unsigned(reg17))}));
              reg73 <= ($signed($signed($signed($unsigned(reg22)))) ?
                  (|(reg65 < $unsigned((reg65 ? reg32 : reg8)))) : (reg24 ?
                      ((|reg8) ^~ $unsigned({(8'hae),
                          wire36})) : ({$unsigned(wire0),
                          (reg55 ^~ reg13)} | $unsigned($unsigned(reg43)))));
              reg74 <= (wire2 ?
                  (^(((reg64 > reg40) < $signed(reg25)) ?
                      wire1 : (reg48 ^ (+reg69)))) : (reg65 >> reg10[(3'h5):(2'h3)]));
            end
          reg75 <= $signed((!$unsigned(reg49[(4'h9):(3'h4)])));
          reg76 <= (|((^{reg73[(4'h8):(1'h1)], $signed(wire2)}) ?
              $unsigned($unsigned($signed(wire4))) : wire0[(1'h1):(1'h0)]));
          if ($unsigned($signed((8'had))))
            begin
              reg77 <= reg58[(2'h3):(2'h2)];
              reg78 <= (^$signed((~|{$unsigned(reg5), reg75})));
              reg79 <= {(+reg19[(1'h1):(1'h0)])};
            end
          else
            begin
              reg77 <= $signed(reg42);
              reg78 <= (~^$unsigned(reg14));
              reg79 <= ((($signed((reg43 | (8'hac))) ~^ reg62) ?
                  (~&{(^wire1),
                      reg62[(5'h16):(4'h8)]}) : (8'ha3)) >> ((((~&reg39) ^~ {reg38,
                      reg31}) ?
                  reg6 : ((^~reg43) ?
                      $unsigned(reg54) : ((8'hb6) ^~ reg67))) && ((-$signed(reg18)) < $unsigned(reg13))));
              reg80 <= $unsigned(reg71[(2'h2):(1'h0)]);
              reg81 <= $unsigned((reg39 ? (8'hb8) : reg62));
            end
          if ($signed($unsigned($signed($signed((~|reg33))))))
            begin
              reg82 <= (reg21[(2'h2):(2'h2)] ?
                  ((7'h48) ?
                      (8'ha5) : $signed(reg10[(3'h5):(3'h4)])) : (reg80 <<< reg13));
              reg83 <= wire3[(1'h1):(1'h0)];
              reg84 <= {(+$signed($signed((!reg17)))),
                  ((reg9[(5'h14):(1'h1)] == $signed((reg27 + reg47))) >>> ($signed($unsigned((8'hba))) >= (^$signed(reg9))))};
            end
          else
            begin
              reg82 <= ((reg67[(4'hb):(2'h2)] ?
                      (($unsigned(reg20) ?
                          $unsigned(reg12) : (reg57 <<< reg37)) && $unsigned(reg5)) : (((reg35 ^~ (8'ha7)) << reg16) ?
                          $unsigned({reg84}) : $unsigned($unsigned(wire4)))) ?
                  reg23[(4'h8):(3'h6)] : reg80[(2'h3):(2'h3)]);
              reg83 <= (~$signed($unsigned((reg14 ?
                  (wire3 ? reg43 : (8'h9e)) : (reg20 ? reg66 : (7'h47))))));
              reg84 <= (reg71[(4'h8):(4'h8)] || $unsigned((&$signed((reg29 ?
                  reg55 : (8'hb0))))));
              reg85 <= ((reg68 ?
                  $unsigned(($signed((8'h9c)) ?
                      reg47[(5'h12):(2'h3)] : reg63[(3'h5):(3'h4)])) : (reg15 | ((8'hac) & {reg57}))) << reg24[(5'h18):(4'hd)]);
            end
        end
      else
        begin
          reg72 <= reg17[(5'h12):(3'h6)];
          reg73 <= reg16[(1'h1):(1'h1)];
          reg74 <= (7'h4c);
          reg75 <= (^reg28[(2'h3):(2'h2)]);
        end
    end
  assign wire86 = {reg39[(3'h4):(2'h3)]};
  always
    @(posedge clk) begin
      if ((((8'hab) || ((~|(reg41 ? (8'haa) : reg13)) ?
          {$unsigned(reg49)} : reg56[(3'h7):(3'h6)])) == reg68[(4'h8):(2'h2)]))
        begin
          reg87 <= $signed(reg32);
          if ((7'h42))
            begin
              reg88 <= ($unsigned(((reg76[(2'h3):(1'h1)] ^~ reg67) <= ({reg52,
                      reg58} ?
                  reg64 : ((8'hbc) ^ reg56)))) + (reg10 ?
                  (((reg51 ?
                      reg30 : wire2) * reg34) || (~(+reg30))) : (~^((+reg13) ?
                      (reg62 | (8'hbe)) : {reg72, reg21}))));
              reg89 <= {((7'h44) ? (8'ha2) : reg80),
                  ($unsigned(((reg13 >>> reg88) > reg41[(4'hf):(3'h6)])) ^ (reg17 + ({(8'hbf),
                      reg60} ^~ {reg83, reg49})))};
            end
          else
            begin
              reg88 <= reg52;
              reg89 <= $unsigned(($unsigned($signed((reg5 != reg67))) ?
                  reg12 : reg60[(4'h9):(3'h4)]));
              reg90 <= {(&(~reg72[(1'h1):(1'h0)]))};
            end
        end
      else
        begin
          reg87 <= (~^$signed($signed(($signed(reg81) >> (reg59 >= reg24)))));
          if (reg47)
            begin
              reg88 <= {reg37[(2'h2):(2'h2)]};
              reg89 <= (reg54[(4'h9):(3'h6)] ?
                  (~(7'h4a)) : reg5[(1'h1):(1'h1)]);
              reg90 <= reg74[(3'h4):(1'h1)];
              reg91 <= $unsigned(reg87[(3'h4):(3'h4)]);
            end
          else
            begin
              reg88 <= $unsigned($signed($signed((8'hb0))));
              reg89 <= $signed(reg72[(2'h3):(2'h3)]);
              reg90 <= $unsigned($unsigned({(reg76 <<< (+reg87)),
                  $unsigned((reg56 >= reg38))}));
              reg91 <= $unsigned((reg70[(1'h0):(1'h0)] ?
                  $unsigned(((reg52 ? (7'h4e) : reg32) || {reg53,
                      (7'h48)})) : ({$unsigned(reg87),
                      (reg41 <<< reg5)} & $signed((reg89 > reg68)))));
            end
          if (($signed((reg63 ^ ($signed((8'ha1)) ?
              {reg60,
                  reg15} : reg55))) << $signed($signed(reg30[(1'h1):(1'h0)]))))
            begin
              reg92 <= (~&reg17[(2'h3):(1'h0)]);
              reg93 <= ($unsigned(($signed((!reg16)) || {reg75[(3'h5):(1'h1)]})) >> $unsigned($signed({reg50,
                  (reg11 ? reg68 : (8'hb9))})));
              reg94 <= $signed(reg20[(4'hf):(4'h9)]);
              reg95 <= {$signed(reg52),
                  (($unsigned(((7'h47) ^ reg73)) & ((reg12 ?
                      reg69 : reg74) >> $unsigned(wire2))) & reg30[(1'h1):(1'h1)])};
            end
          else
            begin
              reg92 <= (^(((wire2 ? reg59 : $unsigned(reg70)) ?
                  reg27[(3'h4):(3'h4)] : $unsigned((~reg19))) || ($signed($unsigned(reg23)) + reg43)));
              reg93 <= $unsigned({$unsigned(reg16),
                  ((^(reg42 ? reg78 : (7'h4b))) ? reg80 : reg40)});
              reg94 <= reg89[(3'h4):(1'h1)];
              reg95 <= (($signed(($unsigned(reg54) - $unsigned(reg94))) >>> reg37) ?
                  $signed((((reg92 | (8'hbe)) || $signed(reg63)) > (~^(reg31 ?
                      reg42 : reg24)))) : {reg76[(3'h7):(1'h1)]});
            end
          if (reg67)
            begin
              reg96 <= (!reg55);
              reg97 <= $unsigned((~|$unsigned((-(|reg11)))));
            end
          else
            begin
              reg96 <= reg42[(3'h6):(3'h6)];
              reg97 <= (!(reg90[(2'h2):(1'h0)] ?
                  ($signed(reg53[(2'h3):(1'h1)]) | reg41) : (|(~|(reg26 || reg70)))));
            end
          reg98 <= $signed(reg49);
          reg99 <= ($unsigned(reg55[(3'h5):(2'h3)]) ?
              ($signed(($signed(reg32) == (reg81 | (8'hbd)))) ?
                  ((((8'hab) ? reg84 : reg35) ?
                          $signed(reg13) : $signed(reg98)) ?
                      (reg93[(1'h1):(1'h0)] ?
                          reg50 : $unsigned(reg16)) : $unsigned(wire3[(2'h3):(1'h1)])) : $signed($unsigned(((7'h46) ?
                      (8'ha0) : reg75)))) : ($unsigned(reg49[(5'h16):(4'he)]) <<< $unsigned($unsigned((reg45 ?
                  reg96 : reg62)))));
        end
      reg100 <= wire3;
      if ((8'hbe))
        begin
          reg101 <= (8'hbd);
        end
      else
        begin
          if ($unsigned(reg68[(4'ha):(4'h8)]))
            begin
              reg101 <= (&($signed(reg58[(2'h2):(1'h1)]) ?
                  $unsigned((+(reg8 ? reg100 : reg62))) : (({reg37, reg40} ?
                      reg83 : (reg93 ? reg74 : reg6)) >= (&reg10))));
              reg102 <= (^reg16[(3'h6):(1'h0)]);
            end
          else
            begin
              reg101 <= reg32[(1'h1):(1'h1)];
              reg102 <= (!$unsigned($unsigned((((8'hbd) ? reg72 : reg73) ?
                  (reg77 >= reg91) : $unsigned((7'h4e))))));
              reg103 <= $signed(((reg22[(3'h6):(3'h5)] ?
                      {reg60[(4'h9):(4'h8)]} : reg26[(1'h1):(1'h0)]) ?
                  (reg27[(3'h7):(3'h7)] ^ $signed({reg67,
                      reg46})) : reg88[(4'hb):(1'h0)]));
              reg104 <= {({$signed((+reg78))} ^ (-(8'hbb)))};
              reg105 <= $signed($unsigned($unsigned($signed(reg82))));
            end
        end
      if (reg54[(4'hd):(3'h7)])
        begin
          if ((~^$unsigned(reg52)))
            begin
              reg106 <= reg6;
              reg107 <= reg84[(3'h5):(2'h3)];
              reg108 <= reg67;
              reg109 <= $unsigned((~|$unsigned($signed(reg14))));
              reg110 <= ($unsigned((($signed(reg88) ?
                      (reg11 <= reg5) : (reg14 ^~ reg64)) < $unsigned($signed(reg40)))) ?
                  ((^~reg50) ?
                      $signed($signed(reg77)) : reg58) : ((^~(reg94[(4'hb):(3'h7)] && (~reg12))) | (^~reg97)));
              reg111 <= reg26;
            end
          else
            begin
              reg106 <= $unsigned(({$signed(reg42),
                  {reg17[(5'h18):(2'h3)], reg82}} <<< $unsigned(reg59)));
              reg107 <= $signed(reg82[(3'h6):(1'h0)]);
            end
          if ($unsigned((((-reg72) ?
                  (((8'hb0) ^ reg73) && reg27[(1'h0):(1'h0)]) : ($signed(reg56) ?
                      $signed((8'hb0)) : (&reg26))) ?
              $unsigned($unsigned((reg43 != reg92))) : {(^~$unsigned(reg61))})))
            begin
              reg112 <= reg20[(4'ha):(2'h2)];
              reg113 <= $signed(({wire1[(1'h0):(1'h0)]} ?
                  ($signed((8'hb9)) ?
                      (8'ha0) : ((reg65 <<< reg110) ?
                          (&reg79) : $signed(reg112))) : {$unsigned($signed(reg6)),
                      (~&(-reg77))}));
              reg114 <= reg46[(5'h10):(4'h8)];
            end
          else
            begin
              reg112 <= {$unsigned(reg55[(3'h7):(3'h5)])};
              reg113 <= ((reg35 ?
                      {((8'ha2) < reg37[(2'h2):(1'h0)])} : $signed(reg79)) ?
                  (7'h45) : $unsigned((~^$signed(reg45))));
              reg114 <= {$unsigned(reg60)};
            end
          reg115 <= $unsigned($unsigned(reg50));
          if ((($signed({reg24[(5'h10):(4'h8)]}) < ((~(reg52 ?
              reg91 : reg64)) <= $signed((reg40 == (7'h41))))) ~^ ((((reg39 ?
                  (7'h4b) : wire3) ?
              (reg60 ?
                  reg115 : reg81) : $unsigned((8'ha1))) <<< $unsigned(reg73)) ^~ (~|($unsigned((8'hb5)) ?
              $unsigned(reg46) : $signed(reg89))))))
            begin
              reg116 <= reg6[(4'ha):(3'h7)];
              reg117 <= $signed(reg102[(4'ha):(4'h8)]);
              reg118 <= ((^(reg114 ?
                  reg65[(4'h8):(2'h2)] : $unsigned(reg20[(2'h2):(1'h1)]))) & (!$unsigned(reg47[(5'h15):(5'h10)])));
              reg119 <= ($unsigned(reg5) ^ reg18[(4'ha):(2'h2)]);
            end
          else
            begin
              reg116 <= (~|$unsigned((&($unsigned(reg103) ?
                  $unsigned(reg13) : (|wire0)))));
              reg117 <= (^~(!(-$unsigned(reg104[(4'he):(4'hb)]))));
              reg118 <= (((({reg90} >= reg68[(3'h4):(2'h3)]) != ({reg106,
                      reg70} ?
                  (+reg26) : (!reg16))) >>> reg22[(2'h3):(2'h2)]) << {($signed(reg87) ?
                      reg51[(4'ha):(3'h4)] : ($signed(reg113) == $unsigned(reg87))),
                  {($signed(reg103) ? (8'hbe) : reg38[(4'hb):(3'h5)])}});
            end
          if ($signed($signed((7'h49))))
            begin
              reg120 <= {$signed($signed((-reg53[(1'h0):(1'h0)])))};
              reg121 <= reg108[(4'hb):(3'h6)];
              reg122 <= $signed((!(((reg99 ?
                      (7'h42) : (7'h41)) >>> $signed(reg19)) ?
                  (reg120[(3'h5):(2'h3)] || reg74) : (!(~|(7'h45))))));
              reg123 <= (wire1 ^ reg70[(2'h2):(1'h1)]);
              reg124 <= ((7'h46) && (|reg54[(5'h11):(5'h10)]));
            end
          else
            begin
              reg120 <= $unsigned(reg54);
            end
          reg125 <= $signed($unsigned(((reg46 || $signed(reg28)) << {$unsigned(reg40),
              $unsigned(reg72)})));
        end
      else
        begin
          if (reg34[(1'h1):(1'h1)])
            begin
              reg106 <= {(~|$unsigned(reg74)),
                  (reg71 >>> (|reg59[(3'h7):(1'h1)]))};
            end
          else
            begin
              reg106 <= {$unsigned(wire1), {$signed(reg35), (8'ha2)}};
              reg107 <= reg28;
              reg108 <= (8'hb3);
            end
          if (((^$signed(reg75)) ?
              (-$unsigned($unsigned((~^reg39)))) : $unsigned($signed($signed((^~reg31))))))
            begin
              reg109 <= reg57;
              reg110 <= $signed(($signed($unsigned(reg15)) <<< reg117[(3'h4):(1'h1)]));
              reg111 <= reg110;
              reg112 <= $signed($signed((wire36[(1'h0):(1'h0)] ?
                  (^~$unsigned(reg51)) : $signed((reg70 ? reg49 : (8'h9e))))));
              reg113 <= $signed((-$signed($unsigned($unsigned(reg56)))));
              reg114 <= reg35;
            end
          else
            begin
              reg109 <= ($signed(($unsigned($signed((8'h9e))) ?
                      {(+(7'h49))} : reg47)) ?
                  (-{reg99[(1'h1):(1'h1)]}) : reg10[(4'hd):(1'h0)]);
              reg110 <= {$signed((($signed(reg20) ^ reg48[(2'h2):(2'h2)]) > ((reg115 - reg66) > $unsigned(reg5))))};
              reg111 <= (|$signed((|$signed($unsigned(reg52)))));
              reg112 <= $unsigned((7'h4e));
            end
        end
      reg126 <= reg113[(3'h4):(1'h1)];
      if (({$signed(((^reg28) ? (reg92 ? reg90 : (8'ha3)) : ((7'h40) - reg79))),
              {$signed(reg59), (reg50 == reg19[(4'hc):(3'h6)])}} ?
          (-(((^reg88) ? (reg45 + reg83) : reg104) ?
              {reg12[(3'h4):(3'h4)]} : $unsigned((7'h44)))) : $signed(reg110[(4'ha):(3'h4)])))
        begin
          if (((~|(~|(^reg60[(3'h7):(3'h4)]))) ?
              (~reg101[(3'h6):(1'h0)]) : reg88))
            begin
              reg127 <= reg19[(3'h4):(3'h4)];
              reg128 <= ($signed(($signed((~&reg105)) ?
                      $unsigned((reg7 ?
                          reg108 : reg80)) : $signed((reg70 & reg78)))) ?
                  $unsigned((|$unsigned((^reg79)))) : (8'ha0));
              reg129 <= $unsigned($signed((reg6 >>> ((~^reg121) ?
                  $signed(reg24) : reg47[(4'hf):(4'hd)]))));
            end
          else
            begin
              reg127 <= {((8'ha6) | (8'h9e)),
                  (wire1 > ((reg85 ?
                      (reg56 ? reg62 : wire3) : (reg18 ?
                          reg47 : reg113)) ~^ reg14))};
              reg128 <= reg16[(2'h2):(2'h2)];
              reg129 <= $unsigned((wire1 < (($unsigned(reg45) >> (8'ha8)) * $unsigned($signed(reg102)))));
              reg130 <= {(reg46[(4'ha):(1'h1)] + reg38),
                  ($signed({(reg128 ? reg67 : reg43)}) ? reg25 : (8'ha6))};
            end
          reg131 <= $unsigned(reg13[(4'ha):(1'h1)]);
        end
      else
        begin
          if ($signed($signed($signed(reg7))))
            begin
              reg127 <= ($unsigned(reg41[(4'h8):(3'h4)]) ~^ $signed({reg47}));
              reg128 <= {$signed((~|$signed(reg122[(5'h10):(4'ha)])))};
              reg129 <= $unsigned($signed($unsigned(reg34)));
              reg130 <= {{{reg32, $unsigned((~reg98))},
                      $unsigned($signed((reg121 ^ reg8)))}};
              reg131 <= ((reg21[(4'hd):(3'h4)] & $unsigned($unsigned($signed(reg35)))) - $unsigned(reg121));
            end
          else
            begin
              reg127 <= wire1[(2'h3):(1'h0)];
              reg128 <= reg62;
              reg129 <= reg94[(3'h7):(3'h6)];
              reg130 <= ((~&($signed($signed(reg118)) ?
                      (~|(|reg42)) : $signed((+reg53)))) ?
                  (&$unsigned(reg25[(4'h9):(3'h4)])) : $signed(($signed($signed(reg15)) ~^ (reg125[(3'h7):(2'h2)] ?
                      reg14 : $signed(reg79)))));
              reg131 <= ((reg53 ^~ $signed($unsigned((wire36 ?
                  reg41 : wire4)))) << reg104[(1'h0):(1'h0)]);
              reg132 <= reg93;
            end
        end
    end
  assign wire133 = reg61[(2'h2):(2'h2)];
  module134 #() modinst939 (.wire138(wire36), .wire137(reg43), .clk(clk), .y(wire938), .wire136(reg35), .wire135(reg103));
  always
    @(posedge clk) begin
      if ((8'hb1))
        begin
          reg940 <= $unsigned($unsigned($unsigned((8'hb4))));
          reg941 <= reg119;
          reg942 <= ({$signed($signed({reg21}))} >= reg941);
          reg943 <= reg77;
        end
      else
        begin
          if (reg132)
            begin
              reg940 <= ((~|reg58) ?
                  $unsigned((($unsigned(reg44) && reg110) && (-reg44[(4'hb):(1'h0)]))) : reg42[(4'ha):(1'h1)]);
            end
          else
            begin
              reg940 <= ($unsigned((~&(8'hbc))) ?
                  ($unsigned((-(reg126 ? reg24 : reg16))) ?
                      $unsigned({(reg32 || reg943),
                          $unsigned(reg18)}) : reg125[(4'he):(4'h8)]) : $unsigned(($unsigned($unsigned(reg131)) > reg25)));
            end
          reg941 <= reg121[(5'h10):(4'hd)];
          if ({$signed((^((8'hb9) ? (^reg20) : reg28))),
              {((~&$signed(reg35)) ?
                      ({reg41,
                          reg73} >> (reg79 <<< (8'ha9))) : $unsigned((reg127 <= reg82))),
                  reg88[(3'h4):(1'h1)]}})
            begin
              reg942 <= ($unsigned((+reg9)) > (reg103 | ($unsigned((+reg940)) ?
                  $unsigned($unsigned(reg102)) : (+reg57))));
            end
          else
            begin
              reg942 <= reg85[(4'hd):(1'h1)];
            end
          reg943 <= ((~|$signed(((8'ha7) ?
              $signed(reg62) : $signed(wire4)))) >> $signed((|($unsigned((7'h4a)) * (8'ha4)))));
        end
      reg944 <= $unsigned(((|reg116) ^~ wire133[(2'h2):(1'h1)]));
      if ((8'hbf))
        begin
          if ((((7'h40) ?
                  $signed(reg124[(4'hc):(4'ha)]) : ($signed((reg60 ?
                          reg124 : reg113)) ?
                      ((~reg24) ~^ {reg15}) : {$signed(reg79)})) ?
              $unsigned((reg85[(3'h7):(1'h1)] <<< wire133)) : {(~($unsigned(reg104) ?
                      (reg130 != reg92) : $unsigned(reg64))),
                  ((^~(+reg90)) ?
                      (reg120[(3'h7):(3'h7)] & (+reg70)) : reg43[(5'h16):(5'h14)])}))
            begin
              reg945 <= $signed({(reg39 >= {(~|reg18),
                      (reg107 ? reg941 : reg51)}),
                  ((^(reg31 ? reg27 : reg41)) <<< reg65)});
              reg946 <= $signed(reg100);
            end
          else
            begin
              reg945 <= (~^($unsigned($signed($unsigned((8'ha0)))) >>> reg123));
              reg946 <= (reg19[(3'h4):(2'h3)] ?
                  (reg93 + $unsigned({$signed(reg121),
                      (reg94 ? reg940 : reg75)})) : $signed(reg111));
            end
          if (reg25[(3'h4):(3'h4)])
            begin
              reg947 <= ((^~((~(wire133 ?
                      reg941 : reg98)) | reg46[(3'h4):(1'h0)])) ?
                  (|reg945[(2'h3):(1'h0)]) : $signed(reg85[(5'h15):(4'hf)]));
              reg948 <= $unsigned(((reg76 ? (^~$signed((8'h9c))) : reg943) ?
                  $unsigned({reg92[(3'h5):(2'h2)],
                      reg110}) : (^($signed(reg44) <<< reg68))));
              reg949 <= ($unsigned($unsigned((|reg8))) | $unsigned((reg55 ?
                  ($unsigned((8'hb1)) >>> (8'ha8)) : reg81)));
            end
          else
            begin
              reg947 <= $signed($signed($signed((+$signed(reg62)))));
              reg948 <= reg77[(5'h18):(4'he)];
              reg949 <= $signed((($signed({reg117}) ^~ (((8'ha8) ?
                      reg16 : reg20) <<< $unsigned(wire36))) ?
                  (8'haf) : (-reg102)));
              reg950 <= $unsigned((($unsigned((reg940 << reg124)) ?
                      $signed({reg27}) : $signed((reg35 ? reg68 : reg49))) ?
                  ({(~&(8'ha4)), (reg94 ? reg68 : reg44)} ?
                      {(~^(8'hab)),
                          (reg33 ?
                              reg96 : reg105)} : reg50) : $unsigned((-reg114[(5'h10):(4'hb)]))));
            end
        end
      else
        begin
          reg945 <= ($signed($unsigned(((reg40 ? reg68 : wire86) <= (wire133 ?
              reg65 : (8'ha2))))) && (reg62 ?
              (7'h40) : (!$unsigned($unsigned(reg105)))));
          reg946 <= ((-reg120[(4'hb):(4'h9)]) ?
              ($signed({$signed((8'ha2))}) >> (~|reg79)) : reg52[(2'h2):(1'h0)]);
          reg947 <= reg7[(4'h8):(2'h3)];
        end
      if ((-reg85[(5'h11):(5'h11)]))
        begin
          if (((~&((reg40 ? (+reg35) : reg89[(1'h1):(1'h1)]) <= reg89)) ?
              ($unsigned($unsigned({reg89})) ?
                  ($signed($signed((7'h49))) ?
                      $signed(reg75) : {(reg22 ? reg73 : wire133),
                          $signed(reg54)}) : (8'hac)) : $unsigned((-reg81))))
            begin
              reg951 <= ((-(-reg78)) < (($signed(reg60[(5'h14):(5'h13)]) ^~ $signed(reg53)) ?
                  ($unsigned((+reg109)) | ((reg10 ~^ reg5) ?
                      (reg72 | (8'hb2)) : $unsigned(reg94))) : reg23[(2'h2):(1'h0)]));
              reg952 <= reg50[(5'h12):(3'h5)];
            end
          else
            begin
              reg951 <= wire4[(1'h1):(1'h1)];
            end
          reg953 <= (~&$unsigned($unsigned(((reg78 ? reg21 : reg948) ?
              reg15[(2'h3):(2'h2)] : reg8))));
          if ($unsigned(reg952))
            begin
              reg954 <= (8'h9c);
              reg955 <= reg81[(4'hd):(4'h8)];
              reg956 <= (~&reg90[(4'ha):(2'h3)]);
              reg957 <= reg131[(4'hf):(2'h2)];
            end
          else
            begin
              reg954 <= (($unsigned($unsigned($unsigned(wire36))) ?
                      $signed($unsigned(reg72[(1'h0):(1'h0)])) : (~reg10[(3'h6):(3'h6)])) ?
                  (reg62 ?
                      (~&$signed(((8'hb2) ?
                          reg38 : reg119))) : $unsigned($unsigned($signed(reg32)))) : ($signed((~(reg952 ?
                      reg71 : reg949))) > ($unsigned((reg75 ?
                      reg62 : reg24)) < (!$unsigned(reg82)))));
              reg955 <= ((((reg69 ?
                      reg127[(3'h6):(2'h2)] : (+wire938)) >= $signed($unsigned(reg53))) ?
                  (~((reg69 ? (7'h48) : reg943) ?
                      (-reg130) : (reg81 ? reg951 : reg63))) : (~^((reg955 ?
                          reg103 : reg24) ?
                      (reg10 ? reg23 : (8'ha2)) : (reg22 ?
                          reg64 : reg17)))) << ((~$unsigned((~&reg9))) ?
                  (&($unsigned(reg83) - (reg13 ?
                      reg82 : reg66))) : reg948[(2'h3):(1'h0)]));
            end
          if (($signed($signed({reg50[(5'h13):(1'h0)]})) > reg54))
            begin
              reg958 <= (8'ha5);
            end
          else
            begin
              reg958 <= (~|$unsigned($unsigned((reg945[(5'h15):(4'hd)] ?
                  $unsigned(reg72) : $signed(reg103)))));
              reg959 <= (reg14[(4'hb):(2'h3)] ?
                  $signed(reg74) : reg124[(5'h12):(3'h5)]);
              reg960 <= reg15[(1'h0):(1'h0)];
            end
          if (reg32)
            begin
              reg961 <= $unsigned(({(wire938 ? reg78 : wire1[(1'h0):(1'h0)]),
                  (reg960[(5'h11):(4'he)] < (reg30 >>> wire36))} << ($signed(((7'h41) || reg25)) ~^ $signed($unsigned(reg31)))));
              reg962 <= (~^$signed((((reg11 ? (8'hac) : reg958) ?
                  reg73[(1'h1):(1'h0)] : $unsigned(reg67)) <<< ((reg11 ~^ reg50) - reg113[(4'h9):(3'h7)]))));
              reg963 <= (reg960 != (^~(((reg958 ? reg99 : (7'h40)) ?
                  (reg69 ?
                      reg60 : reg72) : (~(8'hb3))) && $signed($unsigned(reg113)))));
              reg964 <= ($signed($unsigned(reg34[(5'h13):(4'he)])) ?
                  (({reg37, (^~reg62)} ?
                          $signed((8'haa)) : ($signed((8'ha6)) | (~&reg55))) ?
                      ($unsigned(reg60[(4'hf):(4'h9)]) ?
                          reg110 : reg15[(2'h2):(1'h1)]) : $unsigned((8'hb2))) : reg81[(3'h4):(1'h1)]);
            end
          else
            begin
              reg961 <= $unsigned((^~reg120));
              reg962 <= ((reg117 ?
                      (reg113 ?
                          (&(reg97 ? reg11 : (8'h9d))) : $signed((reg40 ?
                              (7'h44) : reg24))) : $signed($signed($signed((8'h9c))))) ?
                  (8'hb9) : reg10);
              reg963 <= reg124[(4'hd):(4'h8)];
            end
          if ($unsigned($signed((!(|reg126)))))
            begin
              reg965 <= reg958[(3'h5):(1'h0)];
              reg966 <= ($signed({(~^(reg94 ?
                      reg118 : (8'ha8)))}) << (+$unsigned(($unsigned(reg48) ?
                  $signed(reg951) : $unsigned(reg26)))));
              reg967 <= ($unsigned(($unsigned((reg21 ?
                      reg120 : reg19)) | $unsigned((reg114 >> (8'hb0))))) ?
                  $unsigned((((8'h9c) ^~ (^~reg129)) ~^ ({reg46} != (reg27 ?
                      reg44 : reg56)))) : wire3[(1'h0):(1'h0)]);
              reg968 <= reg49[(2'h3):(1'h0)];
              reg969 <= (($signed(reg125) ?
                      $unsigned(reg965[(2'h3):(2'h3)]) : $unsigned((reg961[(2'h2):(2'h2)] ?
                          $signed((8'haf)) : (~&(8'ha1))))) ?
                  reg955[(1'h0):(1'h0)] : reg945);
              reg970 <= $signed(reg80[(4'hd):(4'hc)]);
            end
          else
            begin
              reg965 <= ($unsigned(((~&(reg45 <<< reg970)) == $signed(reg970))) ?
                  $unsigned(wire36) : $signed((($unsigned(reg51) ?
                          (reg940 < reg74) : $signed(reg959)) ?
                      (|reg960) : {(~|reg114), (7'h40)})));
              reg966 <= (reg14[(4'hb):(3'h4)] ?
                  ((!$signed((~^reg72))) + (&(~reg958))) : reg120);
              reg967 <= $unsigned($signed($signed({(7'h4a)})));
              reg968 <= reg113[(4'ha):(3'h6)];
              reg969 <= reg967;
            end
        end
      else
        begin
          reg951 <= reg131;
          reg952 <= reg64;
          if (reg120[(4'h9):(3'h6)])
            begin
              reg953 <= (reg20 ~^ reg120);
              reg954 <= $unsigned(reg942[(4'hc):(3'h7)]);
              reg955 <= $signed($unsigned(reg72));
              reg956 <= {reg945};
            end
          else
            begin
              reg953 <= reg951;
              reg954 <= $signed(reg35[(1'h1):(1'h1)]);
              reg955 <= $unsigned((reg940[(1'h1):(1'h0)] && $signed((~&reg92))));
              reg956 <= ($signed(reg11[(2'h2):(2'h2)]) ?
                  (8'hb2) : $signed($signed($unsigned((reg73 ?
                      reg6 : reg111)))));
              reg957 <= ($signed((reg22 << reg27)) ?
                  reg30 : (reg109[(5'h12):(3'h7)] + (^(^~(+reg37)))));
              reg958 <= (reg966 ?
                  (reg118 <<< reg958) : (&{reg45, reg7[(5'h15):(3'h4)]}));
            end
          reg959 <= $signed({({reg77, (reg959 ? reg95 : reg46)} ?
                  {(&reg53)} : reg100),
              reg110});
          if ((reg947[(4'hb):(3'h4)] && $unsigned((&$signed($unsigned(reg25))))))
            begin
              reg960 <= (reg69[(4'h9):(4'h9)] ? reg94[(3'h4):(2'h2)] : reg55);
              reg961 <= ($signed(({wire4[(1'h1):(1'h1)],
                  {reg97}} ^~ ((reg113 <<< reg103) < (wire938 < reg967)))) > (~(~|reg92)));
              reg962 <= {($signed($signed($signed(reg101))) ?
                      $unsigned($unsigned((reg959 && reg132))) : (reg54 ?
                          reg948 : $unsigned((reg94 ? reg18 : reg956)))),
                  $signed(($unsigned((~&(7'h42))) ?
                      $unsigned((reg29 >= (8'ha9))) : ((~|reg7) - (reg65 ?
                          reg28 : reg60))))};
              reg963 <= {(~(|reg100[(3'h6):(2'h2)]))};
              reg964 <= $signed({(8'hab), $signed(reg43[(1'h0):(1'h0)])});
              reg965 <= reg6[(4'ha):(1'h0)];
            end
          else
            begin
              reg960 <= $signed(($unsigned(reg22[(1'h1):(1'h1)]) >>> reg12[(1'h0):(1'h0)]));
            end
        end
      reg971 <= $signed(reg63[(2'h2):(2'h2)]);
      if (reg23)
        begin
          reg972 <= reg43[(4'hb):(4'hb)];
        end
      else
        begin
          reg972 <= reg112;
          if ($unsigned(reg49[(4'h9):(1'h0)]))
            begin
              reg973 <= (reg75[(3'h5):(1'h1)] == reg121[(3'h6):(3'h6)]);
              reg974 <= ((!(((reg122 <= reg107) ?
                      (~^reg130) : $signed((7'h49))) ?
                  ($signed(reg61) ?
                      reg73 : reg968[(3'h7):(2'h3)]) : {(reg23 | reg951)})) ^ reg48[(4'he):(1'h0)]);
            end
          else
            begin
              reg973 <= $signed(($unsigned(reg52[(1'h0):(1'h0)]) << wire133[(1'h0):(1'h0)]));
              reg974 <= (|(8'hb4));
              reg975 <= ($unsigned(reg59) ?
                  ({reg20} ?
                      $unsigned($signed((~reg75))) : (reg952 ?
                          reg969 : (~^$signed((8'hb9))))) : wire4[(4'ha):(4'ha)]);
              reg976 <= (reg967[(3'h4):(2'h2)] ?
                  reg6[(4'hc):(1'h1)] : {((!reg53) ^ $signed((7'h46))),
                      ($unsigned((reg35 * reg973)) ^ (^{reg58, reg950}))});
              reg977 <= $signed(reg45);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module134
#(parameter param937 = ((~^(((7'h44) ? ((8'haa) != (7'h4d)) : (8'ha3)) >> (~|((8'had) ? (7'h43) : (7'h4e))))) ? (|((((8'hb7) - (8'ha3)) ~^ ((7'h4a) <= (8'hbc))) ? (((8'hab) >= (7'h48)) ? {(8'hbe)} : ((8'h9c) ? (8'hb8) : (8'ha9))) : ((~&(8'hac)) ? ((8'ha0) >= (8'hbe)) : {(8'ha8), (7'h41)}))) : {{({(7'h46)} >= (|(8'ha0))), ((&(8'hbe)) ? ((7'h49) == (8'hac)) : (^~(8'ha0)))}, ((~|{(8'hae)}) ? (((8'haa) | (7'h49)) && ((7'h46) * (8'ha5))) : ({(8'hab)} << {(8'hbb), (8'h9c)}))}))
(y, clk, wire138, wire137, wire136, wire135);
  output wire [(32'h80b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire138;
  input wire [(5'h17):(1'h0)] wire137;
  input wire [(2'h2):(1'h0)] wire136;
  input wire signed [(5'h16):(1'h0)] wire135;
  wire [(5'h1a):(1'h0)] wire936;
  wire signed [(5'h1a):(1'h0)] wire935;
  wire [(5'h1a):(1'h0)] wire925;
  wire signed [(4'hb):(1'h0)] wire924;
  wire [(5'h10):(1'h0)] wire923;
  wire signed [(5'h1a):(1'h0)] wire922;
  wire [(2'h3):(1'h0)] wire913;
  wire [(5'h10):(1'h0)] wire911;
  wire [(4'hd):(1'h0)] wire910;
  wire [(3'h6):(1'h0)] wire909;
  wire signed [(4'ha):(1'h0)] wire907;
  wire [(5'h19):(1'h0)] wire837;
  wire signed [(4'hf):(1'h0)] wire836;
  wire signed [(5'h15):(1'h0)] wire835;
  wire [(4'he):(1'h0)] wire833;
  wire [(5'h14):(1'h0)] wire637;
  wire signed [(4'h9):(1'h0)] wire636;
  wire [(4'hb):(1'h0)] wire197;
  wire signed [(5'h1a):(1'h0)] wire140;
  wire [(4'hf):(1'h0)] wire139;
  wire signed [(3'h7):(1'h0)] wire471;
  wire [(4'ha):(1'h0)] wire473;
  wire signed [(4'hc):(1'h0)] wire634;
  reg [(2'h2):(1'h0)] reg934 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg933 = (1'h0);
  reg [(4'he):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg931 = (1'h0);
  reg signed [(4'he):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg929 = (1'h0);
  reg [(3'h6):(1'h0)] reg928 = (1'h0);
  reg [(4'hb):(1'h0)] reg927 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg926 = (1'h0);
  reg [(4'ha):(1'h0)] reg921 = (1'h0);
  reg [(5'h1a):(1'h0)] reg920 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg919 = (1'h0);
  reg [(2'h3):(1'h0)] reg918 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg915 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg185 = (1'h0);
  reg [(5'h11):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg183 = (1'h0);
  reg [(5'h1a):(1'h0)] reg182 = (1'h0);
  reg signed [(4'he):(1'h0)] reg181 = (1'h0);
  reg [(4'h8):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg177 = (1'h0);
  reg [(5'h10):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg175 = (1'h0);
  reg [(4'h8):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg173 = (1'h0);
  reg [(3'h4):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg170 = (1'h0);
  reg [(5'h10):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg168 = (1'h0);
  reg [(5'h16):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg [(4'ha):(1'h0)] reg165 = (1'h0);
  reg [(3'h7):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg163 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg162 = (1'h0);
  reg [(5'h17):(1'h0)] reg161 = (1'h0);
  reg [(5'h17):(1'h0)] reg160 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg159 = (1'h0);
  reg [(5'h16):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg156 = (1'h0);
  reg [(5'h15):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg154 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg153 = (1'h0);
  reg [(5'h11):(1'h0)] reg152 = (1'h0);
  reg [(5'h17):(1'h0)] reg151 = (1'h0);
  reg [(3'h4):(1'h0)] reg150 = (1'h0);
  reg [(3'h6):(1'h0)] reg149 = (1'h0);
  reg [(3'h4):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg147 = (1'h0);
  reg [(5'h10):(1'h0)] reg146 = (1'h0);
  reg [(2'h2):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg142 = (1'h0);
  reg [(4'hc):(1'h0)] reg141 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg638 = (1'h0);
  reg [(5'h16):(1'h0)] reg639 = (1'h0);
  reg [(5'h15):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg641 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg643 = (1'h0);
  reg [(4'he):(1'h0)] reg644 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg645 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg646 = (1'h0);
  reg [(5'h14):(1'h0)] reg647 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg648 = (1'h0);
  reg [(5'h16):(1'h0)] reg649 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg650 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg651 = (1'h0);
  reg [(4'h9):(1'h0)] reg652 = (1'h0);
  reg [(5'h18):(1'h0)] reg653 = (1'h0);
  reg [(5'h1a):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg656 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg658 = (1'h0);
  reg [(4'hb):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg660 = (1'h0);
  reg [(3'h4):(1'h0)] reg661 = (1'h0);
  reg [(4'h9):(1'h0)] reg662 = (1'h0);
  reg [(4'hc):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg664 = (1'h0);
  reg [(4'he):(1'h0)] reg665 = (1'h0);
  reg [(3'h4):(1'h0)] reg666 = (1'h0);
  reg [(5'h10):(1'h0)] reg667 = (1'h0);
  reg [(5'h17):(1'h0)] reg668 = (1'h0);
  reg [(3'h6):(1'h0)] reg669 = (1'h0);
  reg [(5'h12):(1'h0)] reg670 = (1'h0);
  reg [(3'h6):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg672 = (1'h0);
  reg [(3'h7):(1'h0)] reg673 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg674 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg675 = (1'h0);
  reg [(2'h3):(1'h0)] reg676 = (1'h0);
  reg [(2'h3):(1'h0)] reg677 = (1'h0);
  reg [(5'h12):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg679 = (1'h0);
  reg [(5'h16):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg682 = (1'h0);
  reg [(3'h6):(1'h0)] reg683 = (1'h0);
  reg [(5'h16):(1'h0)] reg684 = (1'h0);
  reg [(4'h9):(1'h0)] reg685 = (1'h0);
  reg [(5'h17):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg687 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg688 = (1'h0);
  assign y = {wire936,
                 wire935,
                 wire925,
                 wire924,
                 wire923,
                 wire922,
                 wire913,
                 wire911,
                 wire910,
                 wire909,
                 wire907,
                 wire837,
                 wire836,
                 wire835,
                 wire833,
                 wire637,
                 wire636,
                 wire197,
                 wire140,
                 wire139,
                 wire471,
                 wire473,
                 wire634,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 reg914,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg638,
                 reg639,
                 reg640,
                 reg641,
                 reg642,
                 reg643,
                 reg644,
                 reg645,
                 reg646,
                 reg647,
                 reg648,
                 reg649,
                 reg650,
                 reg651,
                 reg652,
                 reg653,
                 reg654,
                 reg655,
                 reg656,
                 reg657,
                 reg658,
                 reg659,
                 reg660,
                 reg661,
                 reg662,
                 reg663,
                 reg664,
                 reg665,
                 reg666,
                 reg667,
                 reg668,
                 reg669,
                 reg670,
                 reg671,
                 reg672,
                 reg673,
                 reg674,
                 reg675,
                 reg676,
                 reg677,
                 reg678,
                 reg679,
                 reg680,
                 reg681,
                 reg682,
                 reg683,
                 reg684,
                 reg685,
                 reg686,
                 reg687,
                 reg688,
                 (1'h0)};
  assign wire139 = ((8'h9f) ?
                       (($signed((~^wire136)) == wire138[(3'h4):(2'h3)]) >>> ((~&wire136[(2'h2):(1'h1)]) ?
                           (^wire138) : ((~wire136) >> (wire137 | wire138)))) : {($signed($unsigned(wire136)) >>> {wire138[(3'h6):(1'h0)],
                               {wire136, wire136}})});
  assign wire140 = $signed($signed(((wire139[(4'h9):(3'h7)] && wire138[(2'h2):(2'h2)]) == ((wire138 ?
                           wire137 : wire137) ?
                       (8'hb5) : wire139[(2'h2):(2'h2)]))));
  always
    @(posedge clk) begin
      if ((+($unsigned(($signed(wire137) & wire135[(5'h11):(4'h8)])) ?
          wire138[(4'h8):(2'h2)] : (($unsigned(wire140) <<< (wire138 ?
              wire140 : wire136)) | $signed((wire138 <<< (8'ha3)))))))
        begin
          if (((~|($unsigned(wire140) ?
              ((wire135 || wire135) ?
                  (+wire135) : wire139[(4'ha):(1'h0)]) : $unsigned($unsigned((8'hb3))))) <<< $unsigned($signed($unsigned($unsigned(wire140))))))
            begin
              reg141 <= (!$signed(($signed($signed((7'h4b))) < ((wire138 ^ wire138) - wire136))));
              reg142 <= $signed((wire137[(4'ha):(3'h5)] || (wire135[(1'h1):(1'h0)] ?
                  (!(8'hae)) : ($signed(wire139) >= wire139[(4'he):(3'h6)]))));
              reg143 <= reg142;
              reg144 <= (~&($unsigned(reg142) ?
                  $unsigned(wire135[(4'ha):(2'h3)]) : $signed(wire137)));
            end
          else
            begin
              reg141 <= $unsigned($signed((($signed(wire135) ?
                      (wire136 ? reg141 : reg141) : ((7'h47) == reg142)) ?
                  (wire137 ? (^~reg142) : wire140) : reg141)));
              reg142 <= $signed(($signed((reg141 ?
                  (~^reg142) : $signed(wire139))) | {({reg143,
                      wire140} >>> (wire139 ? wire139 : wire140))}));
              reg143 <= $unsigned($signed(($unsigned((8'ha5)) == wire137[(5'h12):(1'h0)])));
              reg144 <= reg144[(3'h6):(1'h1)];
              reg145 <= ($signed(reg141) ?
                  (reg141[(3'h4):(1'h1)] ?
                      (wire139 ?
                          {wire137[(5'h12):(3'h4)],
                              reg144} : reg141) : ($unsigned((wire139 ?
                              reg142 : reg143)) ?
                          $signed((~wire135)) : wire140)) : wire138);
              reg146 <= (~reg141[(3'h6):(2'h2)]);
            end
        end
      else
        begin
          if (({(8'ha4)} != $signed((8'ha9))))
            begin
              reg141 <= (+reg143);
            end
          else
            begin
              reg141 <= (reg146 != (^~$unsigned($signed($signed(reg143)))));
              reg142 <= reg145;
              reg143 <= $signed(reg142);
              reg144 <= $signed((($unsigned($unsigned(reg143)) >>> (8'hb1)) ?
                  {{(reg143 - reg143)},
                      ($unsigned(wire135) ?
                          $unsigned(reg143) : (wire135 ?
                              wire135 : wire137))} : $unsigned($unsigned(wire135))));
            end
          if ($signed(reg142))
            begin
              reg145 <= reg146[(1'h1):(1'h0)];
              reg146 <= (~^$unsigned((+wire135)));
              reg147 <= (|$signed($signed((wire139 ?
                  {wire136} : $signed(reg142)))));
            end
          else
            begin
              reg145 <= $unsigned((($unsigned((reg145 < (8'hbb))) & (^~(|reg144))) >> $signed(wire138[(3'h4):(1'h0)])));
              reg146 <= wire140;
              reg147 <= reg141[(3'h7):(3'h4)];
              reg148 <= ($signed((|((reg142 ? wire140 : reg143) <<< (wire140 ?
                      reg141 : wire136)))) ?
                  ((reg143[(2'h3):(1'h0)] <= (&wire138)) || $unsigned(wire138)) : $unsigned($unsigned((^~(reg145 ?
                      (7'h47) : reg145)))));
              reg149 <= (|(~(8'haf)));
            end
          reg150 <= ((reg149[(3'h6):(3'h6)] ? reg142[(4'hf):(4'h9)] : (8'h9e)) ?
              $signed(({(wire135 ^ reg141),
                  (+wire140)} || wire140[(5'h14):(5'h14)])) : $unsigned({reg142}));
          if (reg143)
            begin
              reg151 <= $unsigned({$signed((|$signed(reg141)))});
              reg152 <= (reg143 ? $unsigned(reg144[(3'h4):(2'h3)]) : reg144);
              reg153 <= ({(~&(reg145[(2'h2):(1'h0)] >> (~|reg144))),
                      (((wire138 ? reg152 : wire140) ?
                          $unsigned((8'hb5)) : (reg146 + wire137)) >= $signed({wire140}))} ?
                  (($signed((reg145 ^ wire140)) ?
                          $signed(((8'hb2) ?
                              reg147 : wire138)) : $unsigned((8'ha4))) ?
                      ({wire140[(5'h10):(3'h6)],
                          $signed(reg144)} & reg145) : (^~((wire137 || wire136) ?
                          (wire138 ^~ (8'h9f)) : reg150[(1'h0):(1'h0)]))) : (wire138[(3'h4):(3'h4)] ?
                      (!reg147[(3'h7):(1'h1)]) : {(((8'h9c) ?
                              reg143 : reg150) <<< reg143)}));
              reg154 <= (-((~|$signed(((7'h4b) != reg148))) | $unsigned($unsigned((~reg147)))));
              reg155 <= {wire139,
                  {$unsigned(((reg145 + wire135) ?
                          wire138[(3'h4):(1'h1)] : reg150)),
                      (|((8'ha8) ? wire137[(1'h0):(1'h0)] : (~(8'hac))))}};
            end
          else
            begin
              reg151 <= wire136;
            end
          reg156 <= ($signed(reg152[(1'h0):(1'h0)]) ^~ (wire137 - $unsigned($unsigned((~&reg142)))));
        end
      reg157 <= reg145;
      reg158 <= {(($unsigned((reg143 ?
              reg148 : wire137)) < $unsigned($signed(reg148))) <<< $signed({(reg155 - reg142)}))};
      if (reg156)
        begin
          if ($signed($signed(reg155[(4'ha):(3'h6)])))
            begin
              reg159 <= $signed(({(+reg154)} <<< {reg148[(3'h4):(1'h0)]}));
              reg160 <= {((($unsigned(wire138) ^ wire135[(4'he):(4'hc)]) + ((reg150 ?
                              reg145 : wire135) ?
                          (|reg153) : ((8'ha0) ? wire137 : wire138))) ?
                      $unsigned(((8'h9f) * (^~wire136))) : $signed((reg144 | ((7'h4e) ?
                          reg159 : reg147))))};
              reg161 <= (~^(reg152[(4'h9):(2'h3)] & reg146[(1'h1):(1'h1)]));
              reg162 <= {{reg151[(5'h15):(4'hc)],
                      {(reg155[(3'h4):(1'h1)] ?
                              reg159[(2'h2):(1'h0)] : (+reg141)),
                          reg144}}};
            end
          else
            begin
              reg159 <= {$unsigned(wire138)};
            end
        end
      else
        begin
          if ((reg160[(5'h13):(4'he)] ?
              {((wire138 ?
                      (reg150 >>> reg154) : {reg156,
                          reg148}) ^ (+reg143[(1'h1):(1'h1)]))} : (reg153[(1'h0):(1'h0)] ?
                  (~&$unsigned($unsigned(reg146))) : $signed(((reg161 ?
                          wire138 : wire138) ?
                      reg145[(1'h0):(1'h0)] : (~reg141))))))
            begin
              reg159 <= $unsigned(($signed((!(wire138 <= (7'h48)))) ~^ reg156[(2'h3):(1'h1)]));
              reg160 <= (-$signed((reg142[(5'h17):(3'h6)] ?
                  ($unsigned(wire139) ?
                      $signed(wire140) : reg147[(3'h7):(2'h2)]) : (&((8'ha8) ?
                      reg141 : wire137)))));
              reg161 <= (reg153 ? reg143[(1'h1):(1'h1)] : $signed(wire140));
              reg162 <= $signed(((~^((~|(7'h42)) << $signed(reg144))) == ({reg146[(4'hf):(4'h9)],
                  $signed(reg147)} | reg158[(4'hd):(3'h7)])));
              reg163 <= ((wire137 ?
                  (~(8'hb4)) : ({reg142[(5'h12):(2'h3)]} ?
                      reg145 : (^{reg161,
                          reg142}))) <<< (((+$unsigned(reg147)) + reg157[(4'h9):(1'h1)]) ?
                  reg145 : $signed((|wire140))));
            end
          else
            begin
              reg159 <= reg150[(1'h1):(1'h1)];
            end
        end
      if ($unsigned(wire136))
        begin
          reg164 <= $signed(reg149);
          reg165 <= reg153[(3'h7):(2'h3)];
          if ((reg158 - ((((wire138 && reg153) != $signed(reg151)) ?
              ((^~reg158) << (wire139 ?
                  reg146 : reg141)) : ($signed((8'ha0)) & (^~(8'hae)))) <= (reg159 ?
              (~|$unsigned((8'hbe))) : {reg148[(2'h2):(1'h0)],
                  (reg142 ? reg164 : reg163)}))))
            begin
              reg166 <= $unsigned($unsigned({$unsigned($unsigned(reg158))}));
              reg167 <= (reg164[(3'h5):(3'h5)] <<< reg153);
              reg168 <= ((^$unsigned(reg162[(2'h2):(2'h2)])) && ((((+reg143) ?
                      (^~(7'h46)) : (~reg154)) - (~^(~^(8'hb7)))) ?
                  reg155 : $signed((^~$unsigned(reg167)))));
              reg169 <= (&{(((reg168 ? reg162 : wire135) ?
                          reg151 : (reg162 ~^ reg149)) ?
                      reg165[(1'h1):(1'h1)] : ((|reg146) ?
                          $signed(reg161) : (~^wire140)))});
            end
          else
            begin
              reg166 <= wire138;
              reg167 <= $signed($unsigned($signed((reg167[(5'h13):(3'h7)] ?
                  reg154[(4'h8):(3'h6)] : (!wire136)))));
              reg168 <= $signed($unsigned((^(~|$unsigned((7'h42))))));
              reg169 <= ($signed(reg146[(4'hf):(4'ha)]) >= reg144);
              reg170 <= (((reg165 ? {{reg167}, $signed((8'haa))} : (7'h47)) ?
                  reg141 : (^~reg144)) >> ($signed((&reg141)) ?
                  wire137 : reg164[(2'h2):(1'h1)]));
              reg171 <= (-$signed(reg144[(1'h1):(1'h1)]));
            end
          if (wire140)
            begin
              reg172 <= {reg153,
                  ($unsigned($unsigned(reg162[(3'h5):(2'h2)])) ?
                      $unsigned(reg152) : (-reg165))};
              reg173 <= ($signed($unsigned(reg169[(2'h3):(2'h3)])) - reg151);
              reg174 <= $signed((!reg154[(5'h15):(4'hc)]));
              reg175 <= {wire139, reg143[(2'h2):(1'h1)]};
              reg176 <= $signed(($unsigned((^~$unsigned(reg162))) && ({$signed(reg165)} ?
                  $signed(((8'haa) ? reg168 : reg169)) : reg154)));
              reg177 <= reg144[(3'h5):(1'h0)];
            end
          else
            begin
              reg172 <= $signed(reg144);
            end
          if ((8'ha2))
            begin
              reg178 <= $signed(reg150[(1'h0):(1'h0)]);
              reg179 <= (-((($unsigned(reg152) + reg142) ?
                  $signed($signed(reg147)) : (wire135 ?
                      reg171[(4'h9):(4'h8)] : reg162)) | $signed(reg144)));
              reg180 <= $unsigned((reg152[(4'hc):(1'h0)] <<< $unsigned(reg155[(4'hc):(4'hc)])));
            end
          else
            begin
              reg178 <= reg152[(3'h7):(1'h1)];
              reg179 <= (8'hb3);
              reg180 <= (~^$signed($unsigned(reg171)));
            end
        end
      else
        begin
          if (reg146)
            begin
              reg164 <= wire139;
              reg165 <= ($unsigned(reg166[(3'h7):(1'h1)]) ?
                  ({$unsigned($unsigned((7'h43))),
                      {(reg142 == wire140)}} | (reg146[(3'h6):(2'h2)] != (8'hb3))) : (reg162[(4'h8):(4'h8)] ?
                      ($signed(reg165) ?
                          {(reg172 ? (8'hbf) : reg151),
                              wire139} : reg166[(2'h3):(1'h0)]) : reg157[(5'h17):(1'h0)]));
            end
          else
            begin
              reg164 <= (wire135 ^~ (~^$signed($signed({reg163}))));
              reg165 <= $signed(wire140);
              reg166 <= (8'hbf);
              reg167 <= wire136[(1'h1):(1'h1)];
            end
          if ($unsigned(reg169[(2'h3):(2'h2)]))
            begin
              reg168 <= $signed((+reg146[(1'h0):(1'h0)]));
              reg169 <= reg171[(1'h0):(1'h0)];
              reg170 <= $unsigned((^~reg141));
              reg171 <= (+reg146);
              reg172 <= ((~^$unsigned(((8'had) << $signed((8'hb8))))) | ((|reg180) + (~|((8'h9d) >> (8'hb6)))));
            end
          else
            begin
              reg168 <= ((reg146[(3'h4):(2'h3)] ?
                      $signed(($unsigned(reg147) ?
                          reg169 : (reg150 >>> reg171))) : (reg174[(4'h8):(2'h2)] ?
                          $signed($signed(reg174)) : reg149)) ?
                  reg141 : {({$unsigned((7'h46)), (~(7'h49))} ?
                          $unsigned((reg155 ^~ reg174)) : $unsigned((reg176 ?
                              reg157 : reg155)))});
              reg169 <= ((wire140[(5'h16):(4'hc)] ?
                      (reg152[(2'h3):(1'h1)] ?
                          (-(&reg170)) : ((~|reg166) || reg167[(1'h0):(1'h0)])) : (reg162[(3'h6):(1'h0)] && (^(reg156 >> reg146)))) ?
                  (~|reg155) : (~|$unsigned({(reg166 ? reg145 : reg162),
                      (~&reg178)})));
              reg170 <= (-$unsigned({$signed(wire137[(2'h2):(1'h1)]),
                  ((-wire139) ? reg163 : reg178)}));
              reg171 <= {($signed(reg147) > reg157),
                  $signed((reg174 & {wire136, reg156[(5'h10):(3'h5)]}))};
            end
          reg173 <= $signed($signed($unsigned($unsigned({reg148}))));
          reg174 <= ($unsigned(($signed((reg160 ? reg176 : reg148)) ^ {wire140,
              (reg152 | wire137)})) <= reg161[(5'h17):(1'h0)]);
        end
      if ($signed($signed($signed((reg153[(4'h8):(1'h1)] & reg146)))))
        begin
          if (($unsigned((($unsigned(reg177) >= $signed((8'ha0))) & ({reg165} < (|reg169)))) + (8'hb0)))
            begin
              reg181 <= reg165[(2'h3):(2'h2)];
              reg182 <= ($unsigned((($signed(reg162) ?
                  reg159[(1'h0):(1'h0)] : $signed(reg151)) >> wire138)) + $signed(({{wire135,
                          reg173},
                      (reg170 < reg157)} ?
                  $signed((wire136 <<< reg177)) : $unsigned((reg151 ?
                      reg164 : reg166)))));
              reg183 <= $unsigned(({reg146} ?
                  $signed(wire139[(1'h1):(1'h0)]) : $unsigned($unsigned(reg157[(5'h16):(1'h1)]))));
              reg184 <= $unsigned(((reg169[(2'h2):(1'h0)] & reg172[(1'h1):(1'h0)]) ~^ {($unsigned(reg183) >= $unsigned(reg162))}));
              reg185 <= $unsigned((&$unsigned(reg146)));
              reg186 <= $unsigned((&reg155));
            end
          else
            begin
              reg181 <= (~&($signed((reg169 ?
                  (reg174 ? reg167 : reg152) : (reg154 ?
                      wire140 : reg150))) * $unsigned($signed((reg162 ?
                  reg143 : reg186)))));
            end
        end
      else
        begin
          reg181 <= ($unsigned($signed(reg142)) ? (reg150 >= reg163) : reg146);
          if ($unsigned((($signed((reg161 << reg164)) ?
              $signed((^~reg154)) : (reg161[(4'hf):(3'h5)] ?
                  {reg151} : (wire137 ? wire136 : reg175))) & wire140)))
            begin
              reg182 <= (reg160 ?
                  reg175[(3'h5):(2'h2)] : $signed($unsigned({wire140[(4'hd):(4'h9)],
                      $signed((7'h4d))})));
              reg183 <= $signed((~$signed((reg176[(1'h1):(1'h0)] >= $signed((8'had))))));
              reg184 <= ({(!{{reg141}, {reg166}})} >= reg150[(2'h3):(2'h3)]);
              reg185 <= {(8'ha8)};
            end
          else
            begin
              reg182 <= reg181[(1'h1):(1'h0)];
              reg183 <= ($signed((reg168[(4'hb):(4'h9)] + (-$signed(reg152)))) ?
                  (~^($unsigned($unsigned(reg151)) * (&(reg174 ?
                      reg165 : reg143)))) : (8'h9f));
              reg184 <= (+(^$signed($signed(reg156))));
              reg185 <= (8'ha0);
            end
        end
    end
  module187 #() modinst198 (.wire191(reg184), .wire190(reg142), .wire188(reg147), .y(wire197), .clk(clk), .wire192(wire140), .wire189(reg159));
  module199 #() modinst472 (wire471, clk, reg175, reg154, reg158, reg176);
  assign wire473 = $signed({$unsigned(reg154[(5'h12):(4'he)])});
  module474 #() modinst635 (.y(wire634), .clk(clk), .wire476(reg144), .wire478(reg178), .wire477(reg169), .wire475(wire135));
  assign wire636 = $unsigned($signed({reg145, $unsigned(reg186)}));
  assign wire637 = {reg143,
                       ((|((7'h4a) ^~ $unsigned(reg182))) ^~ ($signed($unsigned(reg177)) ?
                           $signed((wire137 == reg186)) : reg175[(4'hf):(4'h8)]))};
  always
    @(posedge clk) begin
      if (wire197[(3'h7):(3'h5)])
        begin
          if ($unsigned($signed((((reg180 ?
              (7'h47) : reg152) - $unsigned(wire137)) * ({reg184} ?
              {wire636} : (reg149 ? (7'h49) : reg174))))))
            begin
              reg638 <= $signed($signed((((reg144 ^ wire636) ?
                  $signed(reg173) : $unsigned(reg178)) > reg165)));
              reg639 <= $signed(reg152);
              reg640 <= reg161[(2'h3):(1'h1)];
              reg641 <= reg143;
              reg642 <= reg178[(5'h17):(4'h8)];
            end
          else
            begin
              reg638 <= reg150;
            end
          reg643 <= {$unsigned(($unsigned(wire136[(1'h0):(1'h0)]) ^~ reg165))};
          reg644 <= ((({$signed(reg156)} >> wire138) <<< ({$unsigned(wire139),
              {reg186, wire137}} || {reg166})) <<< (~&((^~$signed(reg641)) ?
              {(7'h4a), $unsigned(reg175)} : (|$unsigned((7'h40))))));
          if ($signed((|$unsigned($unsigned(((8'h9d) && reg178))))))
            begin
              reg645 <= {($signed(($unsigned((8'hbd)) || (reg158 >>> reg142))) == (8'hbd)),
                  reg150};
              reg646 <= (|$signed(wire138));
              reg647 <= (reg174[(4'h8):(4'h8)] ?
                  $unsigned(reg144[(4'hf):(3'h5)]) : (wire139[(4'hc):(2'h3)] ?
                      reg162[(3'h6):(1'h1)] : reg142[(4'hf):(3'h7)]));
              reg648 <= (-reg173);
              reg649 <= ((8'hac) ? (8'h9d) : $signed(reg151[(5'h17):(4'hb)]));
              reg650 <= (8'ha6);
            end
          else
            begin
              reg645 <= reg171[(4'h8):(1'h0)];
            end
          reg651 <= reg153;
        end
      else
        begin
          if ((~&reg160))
            begin
              reg638 <= ((reg154[(4'h8):(3'h7)] ?
                  (-({reg183, reg172} ?
                      reg176[(4'h9):(3'h5)] : (wire471 | reg175))) : (($signed(reg151) ?
                      (reg645 + reg167) : $signed(reg645)) <<< ($unsigned(reg141) > reg185))) >>> $unsigned(({(reg644 ^ wire636)} ?
                  ((~^reg169) << ((8'hb2) ?
                      reg180 : wire473)) : ((wire138 ^~ wire634) ?
                      $signed(reg178) : $signed(reg144)))));
              reg639 <= {reg149, reg174};
              reg640 <= ($unsigned($unsigned((reg171[(3'h6):(3'h6)] ?
                  $unsigned(reg165) : $unsigned(reg647)))) ^ ($signed(((wire473 > reg182) != (reg147 ~^ reg170))) << ((-reg162) ?
                  reg168[(3'h6):(3'h6)] : (+((8'hbc) < reg167)))));
              reg641 <= reg154[(5'h13):(4'hc)];
              reg642 <= $unsigned((+((wire473[(2'h2):(1'h1)] && $signed(reg174)) - ((reg183 << reg162) & (^~reg639)))));
              reg643 <= {($signed(wire140) | {$unsigned($signed(reg149))}),
                  reg165};
            end
          else
            begin
              reg638 <= ((reg150[(2'h3):(1'h0)] > ((!reg169[(3'h6):(3'h4)]) ?
                  ((wire471 ? reg151 : wire637) ?
                      $unsigned(reg638) : (^~reg170)) : ($unsigned(reg650) < (reg170 == reg143)))) && reg154[(5'h15):(5'h11)]);
              reg639 <= {$unsigned(reg181),
                  {(reg645[(2'h2):(1'h1)] ?
                          ({reg647, reg152} ?
                              wire197 : (reg643 ?
                                  reg166 : reg153)) : wire135[(5'h15):(5'h12)]),
                      reg642[(3'h6):(2'h2)]}};
              reg640 <= {(reg158[(1'h1):(1'h0)] ? {{(^wire197)}} : reg172)};
              reg641 <= wire135;
            end
          if ({reg146[(4'ha):(3'h6)]})
            begin
              reg644 <= wire135;
            end
          else
            begin
              reg644 <= reg183[(3'h6):(2'h3)];
              reg645 <= reg171[(4'he):(4'he)];
              reg646 <= $unsigned(($unsigned((^(^~(8'hb0)))) < (~($unsigned((8'h9f)) ?
                  $signed((7'h46)) : reg142[(4'ha):(4'ha)]))));
              reg647 <= (^~({$unsigned((&reg149)),
                  $signed($unsigned(reg156))} << $signed(((reg161 ?
                  reg161 : wire139) | (reg180 | reg171)))));
            end
          if ($signed(reg639))
            begin
              reg648 <= ($unsigned($unsigned($unsigned((^reg146)))) ~^ (7'h43));
            end
          else
            begin
              reg648 <= (reg185[(3'h4):(2'h2)] < reg643);
              reg649 <= wire634[(3'h6):(1'h0)];
              reg650 <= $signed({(reg155[(5'h10):(5'h10)] ^ $signed((&reg175)))});
              reg651 <= reg171;
              reg652 <= (7'h47);
            end
        end
      if ((-(7'h47)))
        begin
          reg653 <= reg141[(3'h5):(2'h3)];
          reg654 <= (~$signed((+reg146)));
          if ((|($unsigned(($unsigned(reg162) ?
                  (wire471 >> reg170) : (reg167 ? reg153 : reg150))) ?
              wire636[(2'h3):(2'h2)] : $signed(reg164))))
            begin
              reg655 <= ($signed($signed({reg166[(2'h3):(1'h1)]})) ?
                  ($signed(wire197) ?
                      $signed((8'hba)) : wire136[(1'h0):(1'h0)]) : ($unsigned((8'ha7)) ?
                      (reg153 << (8'hbb)) : $unsigned(reg165[(2'h2):(1'h1)])));
              reg656 <= (^{(reg146 ?
                      ($unsigned(wire138) <= reg160) : wire636[(2'h2):(1'h1)])});
            end
          else
            begin
              reg655 <= $signed(($unsigned(($unsigned(reg148) <<< (8'ha6))) == ((((7'h4a) ?
                      wire637 : (7'h46)) ?
                  $signed(reg644) : (wire136 ?
                      (8'hbe) : reg162)) != reg144[(4'h8):(2'h3)])));
              reg656 <= $signed($signed(((~&(reg173 & reg156)) >= ($unsigned(reg648) ?
                  reg165[(3'h7):(2'h3)] : $unsigned(reg145)))));
              reg657 <= (~$signed(({reg652,
                  wire140} ~^ $signed($unsigned(reg167)))));
              reg658 <= ($signed($signed(($unsigned(reg168) ?
                  (!(7'h40)) : reg655[(3'h7):(2'h3)]))) == {(~^(^(reg639 && reg161)))});
            end
          if ((((+reg183) ?
                  $unsigned(reg639[(4'hd):(3'h4)]) : {$signed({(7'h4a),
                          reg651}),
                      {reg178}}) ?
              (!((^~wire471[(2'h3):(2'h2)]) ?
                  reg638 : ((^reg171) ?
                      reg167 : (reg155 ?
                          reg639 : (8'ha0))))) : ((~|$unsigned(((8'hbd) ?
                      reg146 : (8'hba)))) ?
                  reg177[(3'h7):(1'h0)] : $signed(reg151))))
            begin
              reg659 <= reg653;
              reg660 <= (8'ha2);
              reg661 <= wire471[(3'h7):(1'h0)];
              reg662 <= wire135[(1'h1):(1'h1)];
              reg663 <= wire140[(4'hf):(4'h8)];
              reg664 <= $unsigned((~&$unsigned(reg644[(3'h4):(2'h3)])));
            end
          else
            begin
              reg659 <= (((~$signed((^reg178))) == (reg171 & reg643)) ?
                  ((reg179 < (~^$signed(reg653))) <= $signed((8'ha9))) : reg141);
              reg660 <= (-{(!$unsigned(reg186[(5'h12):(5'h10)]))});
              reg661 <= $unsigned($unsigned(reg163));
              reg662 <= reg644[(3'h7):(3'h7)];
              reg663 <= ($unsigned($signed(((reg648 ?
                      reg170 : (8'hb5)) & $signed(reg162)))) ?
                  (((^~(reg153 + reg177)) ?
                          $signed((reg651 ? (8'hb7) : reg653)) : ((reg172 ?
                                  reg165 : reg654) ?
                              $signed(reg176) : (reg174 | reg179))) ?
                      $unsigned($signed(((8'h9f) < wire136))) : ((wire140 ?
                          (^~reg649) : reg161[(3'h7):(3'h7)]) - $unsigned($signed(reg172)))) : ((~&{(wire140 >= reg164),
                      (reg153 * wire636)}) << reg650));
              reg664 <= reg174;
            end
          if ($signed((^(+$signed($unsigned((8'ha5)))))))
            begin
              reg665 <= reg642;
              reg666 <= reg177;
            end
          else
            begin
              reg665 <= (((8'ha8) ?
                      reg155[(3'h4):(2'h2)] : (|reg153[(3'h5):(2'h3)])) ?
                  $signed($unsigned((reg169[(4'ha):(2'h2)] <<< $unsigned(reg157)))) : (|(($unsigned(reg148) == (reg170 ?
                      reg152 : reg143)) ^~ reg151[(4'he):(3'h5)])));
              reg666 <= reg174[(3'h5):(2'h3)];
              reg667 <= $unsigned({(!reg174[(1'h0):(1'h0)])});
              reg668 <= {(!{(|((7'h41) - reg186)),
                      ((7'h49) ? $unsigned(reg651) : $signed(wire197))}),
                  (({$signed(reg649),
                      reg148} >= (+(7'h46))) > $signed({reg168[(4'h9):(3'h7)],
                      reg149[(2'h3):(1'h0)]}))};
              reg669 <= $unsigned((~|((reg178[(4'hd):(4'hd)] ?
                      (reg649 ? wire135 : reg156) : $signed(reg175)) ?
                  wire138[(2'h3):(1'h0)] : reg653)));
            end
          if ($signed((!(8'hae))))
            begin
              reg670 <= ((reg162 || wire139) ^~ $signed($signed((&((8'hb6) <= wire636)))));
              reg671 <= (reg175[(3'h6):(3'h6)] ?
                  (~&(~^(~((8'hbf) || wire637)))) : reg650);
            end
          else
            begin
              reg670 <= $signed((((reg171 ?
                  $signed(reg658) : (reg175 ?
                      reg170 : reg146)) ^ wire197[(4'hb):(3'h4)]) >>> reg671));
            end
        end
      else
        begin
          reg653 <= ($signed((($signed((7'h45)) ?
                  $unsigned(reg639) : reg144) ^~ reg154[(4'ha):(2'h2)])) ?
              $unsigned((+((wire634 ? reg647 : reg663) ?
                  (&reg641) : (~(8'ha6))))) : reg159[(1'h0):(1'h0)]);
          if (reg174)
            begin
              reg654 <= reg639;
              reg655 <= {$signed(reg183[(1'h1):(1'h1)]), reg182};
              reg656 <= (reg650 & (^~reg151));
              reg657 <= reg143;
            end
          else
            begin
              reg654 <= wire636[(1'h1):(1'h0)];
            end
          if ($unsigned((^(|reg641[(1'h0):(1'h0)]))))
            begin
              reg658 <= $signed(reg163);
              reg659 <= {($unsigned(($unsigned(reg662) * (reg158 && reg658))) ?
                      reg662 : $signed(reg178[(1'h1):(1'h1)]))};
              reg660 <= ($unsigned(reg656) ~^ (~reg659[(1'h1):(1'h0)]));
              reg661 <= (~&(8'hb7));
            end
          else
            begin
              reg658 <= $signed(($signed((|$signed((8'ha5)))) ?
                  $unsigned(wire473[(2'h3):(2'h2)]) : $signed($signed(reg667))));
            end
          reg662 <= (^~reg666);
          if (reg668)
            begin
              reg663 <= $unsigned(reg160[(1'h1):(1'h1)]);
              reg664 <= ($unsigned(reg665[(4'h8):(1'h0)]) | (~reg150));
              reg665 <= (reg151[(1'h0):(1'h0)] ?
                  reg146[(4'hd):(1'h1)] : reg156[(4'hb):(3'h7)]);
              reg666 <= (8'ha8);
              reg667 <= reg659[(3'h4):(3'h4)];
              reg668 <= $unsigned((~^$unsigned(reg639)));
            end
          else
            begin
              reg663 <= {$unsigned($unsigned(($signed(reg650) >>> {reg671})))};
              reg664 <= (|wire197[(1'h1):(1'h1)]);
              reg665 <= {(wire634 * $unsigned(($signed((8'ha6)) ?
                      (&reg159) : reg173)))};
              reg666 <= reg169[(4'hd):(1'h0)];
              reg667 <= reg646;
            end
          if (reg643)
            begin
              reg669 <= $unsigned((8'hbd));
              reg670 <= (7'h46);
              reg671 <= wire135[(3'h7):(3'h4)];
              reg672 <= $unsigned((!(7'h48)));
            end
          else
            begin
              reg669 <= $unsigned(reg646[(1'h0):(1'h0)]);
              reg670 <= $signed((&(((-reg144) << (~^reg642)) ?
                  $unsigned($signed((7'h42))) : reg175[(4'hf):(1'h0)])));
              reg671 <= {reg168};
              reg672 <= reg162;
              reg673 <= $signed((|$unsigned((reg185[(5'h10):(4'hc)] ?
                  (reg141 ? wire138 : wire471) : reg148[(1'h1):(1'h1)]))));
              reg674 <= (+reg144[(3'h5):(3'h5)]);
            end
        end
      if ({{(reg672[(4'hb):(4'h8)] ?
                  ((reg182 < reg173) ?
                      (wire140 >>> reg665) : (reg656 ?
                          (8'hb8) : reg174)) : reg672),
              wire135}})
        begin
          reg675 <= reg647;
          if ($signed(reg645))
            begin
              reg676 <= reg642[(3'h5):(3'h5)];
              reg677 <= reg167;
            end
          else
            begin
              reg676 <= $signed($signed((7'h44)));
              reg677 <= $unsigned((((&reg666[(2'h2):(1'h1)]) ?
                  ({reg185,
                      reg181} + (reg671 == (8'hb0))) : reg655[(3'h6):(3'h6)]) >> ((~^reg184[(4'hc):(1'h0)]) || $unsigned($unsigned(reg162)))));
              reg678 <= {wire138};
              reg679 <= ($signed(reg156) && $signed(((|$unsigned(reg172)) ?
                  wire135 : (((8'ha6) ? reg655 : reg652) ?
                      (reg676 ? reg159 : wire136) : reg666[(2'h2):(1'h1)]))));
              reg680 <= (reg163[(3'h7):(3'h4)] * reg643);
            end
          if ((reg152 == $unsigned($unsigned(reg173[(5'h15):(2'h3)]))))
            begin
              reg681 <= $unsigned((&$signed(($signed(reg167) != {(7'h42),
                  reg144}))));
              reg682 <= (reg649 ? reg679 : (~&reg646[(2'h3):(2'h2)]));
            end
          else
            begin
              reg681 <= reg145;
            end
          if ((~|(8'hba)))
            begin
              reg683 <= wire471;
              reg684 <= reg141;
              reg685 <= reg662;
              reg686 <= $signed((reg648 ?
                  reg176[(1'h1):(1'h1)] : (~|{$signed(reg638),
                      $unsigned(wire471)})));
              reg687 <= reg142;
              reg688 <= (($signed((reg669[(1'h1):(1'h1)] ?
                  $unsigned(reg173) : reg659[(1'h0):(1'h0)])) == $signed({$unsigned(reg147)})) != (($signed($unsigned((8'ha6))) <= $unsigned((reg686 || reg670))) ?
                  (~^($unsigned(reg166) ?
                      reg663 : (reg160 ? reg647 : reg146))) : reg639));
            end
          else
            begin
              reg683 <= reg665[(4'h9):(2'h2)];
              reg684 <= (|(-reg153));
            end
        end
      else
        begin
          if ((((~&reg147) ?
                  (reg148[(1'h0):(1'h0)] >>> ((&reg172) ?
                      (wire637 ?
                          reg648 : reg180) : $unsigned(reg173))) : ({((8'ha5) != (8'ha5))} ?
                      $signed($signed(reg644)) : (reg652[(3'h7):(2'h3)] & $unsigned(reg672)))) ?
              (($unsigned($unsigned(reg661)) ?
                      reg674[(4'ha):(2'h2)] : ((wire637 - wire634) ?
                          wire137 : {reg667, reg157})) ?
                  ((~|(+wire634)) ?
                      $unsigned({reg150}) : reg661[(2'h3):(1'h0)]) : reg167) : $unsigned(($signed($signed(reg652)) >> ($signed(reg676) >> $signed((8'hb3)))))))
            begin
              reg675 <= (reg656[(5'h10):(4'h9)] ?
                  {(&reg664),
                      $unsigned((~$unsigned(reg145)))} : $unsigned((~|((reg684 && reg679) ?
                      (!reg655) : (wire140 << reg646)))));
              reg676 <= $signed($signed($unsigned(({reg645, reg638} ?
                  {reg665, reg647} : reg176[(2'h2):(1'h1)]))));
            end
          else
            begin
              reg675 <= reg183[(3'h5):(1'h1)];
              reg676 <= reg662;
            end
          reg677 <= $unsigned(reg162);
        end
    end
  module689 #() modinst834 (.clk(clk), .wire692(reg643), .wire694(reg688), .y(wire833), .wire690(reg149), .wire691(reg165), .wire693(reg158));
  assign wire835 = (+($unsigned(reg648[(3'h5):(3'h5)]) ?
                       ((~&reg177[(3'h4):(2'h3)]) ?
                           reg681[(1'h1):(1'h1)] : $signed({reg664})) : $signed($unsigned((7'h45)))));
  assign wire836 = (^$signed(reg661));
  assign wire837 = reg657;
  module838 #() modinst908 (.wire843(reg653), .wire840(reg639), .wire842(reg182), .wire841(reg684), .y(wire907), .wire839(reg664), .clk(clk));
  assign wire909 = (~^({(^~(|reg671))} + {(!{wire137, reg638})}));
  assign wire910 = (&reg667);
  module187 #() modinst912 (wire911, clk, reg163, reg688, reg650, reg687, reg680);
  assign wire913 = (((reg675[(3'h6):(2'h2)] - $signed($signed(reg683))) ^ (&reg172[(1'h0):(1'h0)])) && (|($signed((reg157 - (8'haf))) | (reg650[(5'h11):(4'hd)] > reg170))));
  always
    @(posedge clk) begin
      if ({reg172})
        begin
          reg914 <= reg157;
          if ($unsigned($unsigned(($unsigned((&(8'h9c))) > ((reg662 <<< reg175) ^ (-wire634))))))
            begin
              reg915 <= (^$signed((^{(reg673 >> reg172), reg157})));
              reg916 <= $unsigned(($unsigned((!$unsigned(wire833))) << ($unsigned(wire135) ?
                  $signed((reg152 ? reg169 : reg660)) : ({wire837} >> {(8'hb0),
                      reg668}))));
              reg917 <= $unsigned($signed({$unsigned($signed(reg162))}));
            end
          else
            begin
              reg915 <= (~&reg145[(2'h2):(1'h1)]);
            end
          if ({$unsigned((^$signed({wire139}))), (~{reg176})})
            begin
              reg918 <= $signed(reg180[(2'h3):(2'h2)]);
            end
          else
            begin
              reg918 <= wire473;
              reg919 <= (($unsigned(reg685) == {reg655[(4'hc):(4'hc)]}) ?
                  $unsigned((8'hb5)) : (7'h48));
              reg920 <= ($unsigned({$signed(reg144[(4'hd):(3'h7)]),
                  reg685}) | (reg178 <= wire473[(4'h9):(2'h3)]));
              reg921 <= reg156;
            end
        end
      else
        begin
          reg914 <= (((reg143[(5'h16):(3'h6)] <= ((reg920 ?
                  reg165 : (8'hbc)) >= reg650)) ?
              ((-$signed(reg167)) - ((&reg672) > (+(7'h42)))) : ((~^{wire836,
                  reg914}) != reg165[(2'h2):(1'h1)])) >= $unsigned(reg178));
        end
    end
  assign wire922 = $signed(($signed(reg182[(2'h3):(1'h0)]) >>> $unsigned({((7'h4b) ?
                           reg158 : reg661),
                       $unsigned(reg173)})));
  assign wire923 = wire835;
  assign wire924 = $signed(reg143[(5'h15):(3'h4)]);
  assign wire925 = $unsigned(reg171[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ($unsigned(({reg180[(3'h6):(2'h2)],
          (&(reg668 ^ reg666))} || {(^(wire138 > wire922)), {reg185}})))
        begin
          if (reg145[(2'h2):(1'h1)])
            begin
              reg926 <= ((~|({$signed(reg652), reg173} ?
                  ($signed(wire637) ?
                      (reg662 ?
                          wire637 : reg160) : reg676) : {(reg170 * wire138),
                      $unsigned(wire634)})) >>> (~|($signed(((8'hba) ?
                      wire139 : reg157)) ?
                  $unsigned(reg659[(3'h5):(1'h0)]) : $unsigned((reg649 ?
                      reg186 : reg158)))));
              reg927 <= reg662[(3'h7):(3'h4)];
              reg928 <= $unsigned(({(reg640 ?
                          wire835[(5'h10):(4'hd)] : (8'ha2)),
                      $unsigned((&reg159))} ?
                  ((~(reg675 ? reg921 : reg141)) ?
                      wire835 : (((8'h9d) ?
                          reg669 : reg156) ^~ {wire135})) : (reg676[(1'h1):(1'h1)] ?
                      $signed((reg667 ^~ reg649)) : ((reg661 + wire837) ?
                          reg150[(3'h4):(2'h2)] : reg645))));
              reg929 <= reg165[(1'h1):(1'h1)];
            end
          else
            begin
              reg926 <= ($signed((reg914[(2'h3):(2'h3)] ?
                  ((reg160 ? reg149 : (8'h9f)) ?
                      $signed(reg677) : $unsigned(reg186)) : (reg166[(2'h3):(1'h0)] ?
                      {reg667} : (reg141 ?
                          reg148 : (8'h9c))))) >> reg185[(4'hc):(3'h7)]);
              reg927 <= (reg664 ?
                  ($signed($unsigned($signed(reg921))) ?
                      {(!{(8'hbb)})} : reg177[(4'hb):(1'h1)]) : $signed({(((8'ha9) >>> reg178) ?
                          (wire907 ?
                              reg670 : (7'h4d)) : reg647[(2'h3):(1'h1)])}));
              reg928 <= reg920[(4'h8):(1'h0)];
              reg929 <= (reg656[(1'h0):(1'h0)] ?
                  $signed($signed({reg919,
                      $signed(reg172)})) : reg175[(2'h2):(1'h0)]);
              reg930 <= reg927[(2'h3):(1'h1)];
            end
        end
      else
        begin
          reg926 <= $signed(reg175[(3'h4):(2'h3)]);
          reg927 <= $unsigned($unsigned($unsigned($signed(((8'h9c) <= reg641)))));
          if ((((-(wire471 > (&(8'hb2)))) + reg677) ?
              (+reg678[(1'h1):(1'h0)]) : ($unsigned(((reg657 ?
                  reg645 : reg661) - wire836)) && reg643)))
            begin
              reg928 <= $signed(($unsigned(reg646[(3'h4):(3'h4)]) ?
                  $signed(reg152) : (7'h46)));
              reg929 <= $unsigned($unsigned($unsigned(wire637[(1'h1):(1'h0)])));
              reg930 <= $unsigned(reg157);
              reg931 <= (reg656[(1'h1):(1'h0)] ?
                  reg666 : $unsigned({$signed($unsigned(reg662)),
                      ({wire637, reg161} <= reg653)}));
            end
          else
            begin
              reg928 <= $signed((&((+wire837[(5'h19):(3'h4)]) >>> ((reg667 <= reg683) ?
                  (reg662 ? (7'h48) : (8'hac)) : {reg670}))));
            end
          reg932 <= $unsigned(($unsigned(({reg680, (7'h44)} ?
              (^~reg149) : (-wire923))) == (~|{reg930[(4'h8):(3'h5)]})));
          reg933 <= $unsigned(($signed(($signed(reg152) ^~ (reg665 ^ reg638))) <= wire925));
        end
      reg934 <= ((reg177 ^~ reg646) <<< reg182);
    end
  assign wire935 = reg932[(3'h6):(2'h3)];
  assign wire936 = $signed((((wire833 ? (reg929 << reg175) : (^~reg679)) ?
                           $signed($unsigned(reg157)) : $signed($signed(reg158))) ?
                       ($unsigned((7'h4a)) ?
                           (&reg678[(3'h4):(3'h4)]) : wire833[(2'h2):(2'h2)]) : wire137[(4'h9):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module838  (y, clk, wire843, wire842, wire841, wire840, wire839);
  output wire [(32'h3e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire843;
  input wire signed [(5'h19):(1'h0)] wire842;
  input wire signed [(5'h16):(1'h0)] wire841;
  input wire [(4'hf):(1'h0)] wire840;
  input wire signed [(5'h13):(1'h0)] wire839;
  wire [(3'h6):(1'h0)] wire906;
  wire [(4'ha):(1'h0)] wire864;
  wire [(5'h16):(1'h0)] wire863;
  wire signed [(5'h15):(1'h0)] wire862;
  wire signed [(5'h16):(1'h0)] wire861;
  wire [(4'hb):(1'h0)] wire860;
  wire signed [(5'h10):(1'h0)] wire859;
  wire [(5'h12):(1'h0)] wire858;
  wire signed [(4'hf):(1'h0)] wire857;
  wire signed [(5'h18):(1'h0)] wire856;
  wire [(5'h18):(1'h0)] wire854;
  wire [(4'hd):(1'h0)] wire845;
  wire [(4'h9):(1'h0)] wire844;
  reg [(5'h15):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg902 = (1'h0);
  reg [(5'h11):(1'h0)] reg901 = (1'h0);
  reg [(4'h8):(1'h0)] reg900 = (1'h0);
  reg [(5'h1a):(1'h0)] reg899 = (1'h0);
  reg [(5'h13):(1'h0)] reg898 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg897 = (1'h0);
  reg [(5'h11):(1'h0)] reg896 = (1'h0);
  reg [(5'h19):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg894 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg893 = (1'h0);
  reg [(5'h12):(1'h0)] reg892 = (1'h0);
  reg [(5'h17):(1'h0)] reg891 = (1'h0);
  reg [(5'h11):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg889 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg887 = (1'h0);
  reg [(4'h8):(1'h0)] reg886 = (1'h0);
  reg [(3'h5):(1'h0)] reg885 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg884 = (1'h0);
  reg [(5'h13):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg882 = (1'h0);
  reg [(5'h10):(1'h0)] reg881 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg880 = (1'h0);
  reg [(2'h2):(1'h0)] reg879 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg878 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg876 = (1'h0);
  reg [(3'h6):(1'h0)] reg875 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg874 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg873 = (1'h0);
  reg [(5'h1a):(1'h0)] reg872 = (1'h0);
  reg [(2'h3):(1'h0)] reg871 = (1'h0);
  reg [(5'h12):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg869 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg868 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg867 = (1'h0);
  reg signed [(4'he):(1'h0)] reg866 = (1'h0);
  reg [(5'h1a):(1'h0)] reg865 = (1'h0);
  reg [(3'h7):(1'h0)] reg855 = (1'h0);
  reg [(2'h2):(1'h0)] reg853 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg852 = (1'h0);
  reg [(5'h1a):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg850 = (1'h0);
  reg [(5'h14):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg848 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg847 = (1'h0);
  reg [(3'h6):(1'h0)] reg846 = (1'h0);
  assign y = {wire906,
                 wire864,
                 wire863,
                 wire862,
                 wire861,
                 wire860,
                 wire859,
                 wire858,
                 wire857,
                 wire856,
                 wire854,
                 wire845,
                 wire844,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg855,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 (1'h0)};
  assign wire844 = (&((wire841 ?
                           wire843[(3'h4):(1'h1)] : ({(8'hb0)} ?
                               wire842[(3'h5):(3'h5)] : $signed(wire842))) ?
                       wire843 : $unsigned((|(wire840 + wire839)))));
  assign wire845 = wire844[(4'h9):(2'h3)];
  always
    @(posedge clk) begin
      if ($signed(($signed({(8'hbe)}) ?
          ((wire840[(2'h3):(1'h0)] ? $signed(wire845) : (wire840 != wire843)) ?
              $unsigned(wire842[(1'h0):(1'h0)]) : $unsigned((wire843 >= wire845))) : $signed(wire845[(4'hd):(3'h4)]))))
        begin
          if ($signed(wire844[(4'h8):(1'h1)]))
            begin
              reg846 <= (^(~{(|$signed(wire839))}));
              reg847 <= (|$unsigned((-((~wire844) | (8'ha2)))));
              reg848 <= wire842[(1'h0):(1'h0)];
              reg849 <= $unsigned(reg847[(2'h2):(1'h0)]);
              reg850 <= $signed(wire839[(4'he):(4'h9)]);
              reg851 <= (wire845 ?
                  wire839[(3'h7):(2'h2)] : {(-$signed({wire840, reg850}))});
            end
          else
            begin
              reg846 <= ($unsigned((7'h4b)) < ((+reg847[(2'h2):(2'h2)]) < (wire844[(4'h9):(2'h2)] ?
                  wire845 : (reg849[(4'h9):(2'h3)] + (wire842 + wire844)))));
              reg847 <= {wire844};
              reg848 <= $unsigned({(+wire842[(5'h10):(4'h9)])});
              reg849 <= reg848;
            end
          reg852 <= (7'h4a);
          reg853 <= (~&(8'hb9));
        end
      else
        begin
          if (({(|wire839[(4'hc):(3'h7)])} ?
              (wire844 == (8'hb4)) : $unsigned(reg850)))
            begin
              reg846 <= $signed(($signed(($signed(wire843) ?
                  reg847 : (reg846 < wire839))) && $signed(wire842)));
            end
          else
            begin
              reg846 <= (+{reg850});
              reg847 <= $unsigned((((~&{(8'hbc), reg853}) ?
                      reg853 : reg852[(4'hc):(4'hb)]) ?
                  $unsigned((~^wire843)) : {((7'h4a) <<< (reg846 ^~ wire839)),
                      $unsigned($unsigned(reg846))}));
              reg848 <= $signed($unsigned((wire845[(4'h8):(3'h6)] ?
                  (^~{reg846, reg850}) : wire842[(4'hd):(4'hc)])));
              reg849 <= reg853[(1'h1):(1'h0)];
              reg850 <= (reg847 == reg846[(2'h3):(2'h3)]);
              reg851 <= wire840[(2'h3):(2'h2)];
            end
          reg852 <= {((|reg851) ?
                  wire843[(4'hc):(3'h6)] : (~$signed($signed(wire841))))};
          reg853 <= {$unsigned(($unsigned((wire839 & wire845)) >> $unsigned(reg847[(2'h3):(1'h1)])))};
        end
    end
  assign wire854 = ($unsigned(wire843) <<< $unsigned(reg850));
  always
    @(posedge clk) begin
      reg855 <= wire845;
    end
  assign wire856 = ({($unsigned(wire839) ?
                           (&$signed(reg849)) : $unsigned($unsigned(reg855)))} != $signed((~$unsigned(wire844[(1'h1):(1'h0)]))));
  assign wire857 = $unsigned($unsigned(wire844));
  assign wire858 = $unsigned({$unsigned(((reg853 && reg850) > reg851)),
                       (reg852[(4'ha):(2'h2)] == (~&$signed(reg851)))});
  assign wire859 = $unsigned(($signed(wire845[(2'h2):(1'h1)]) && (-(^(wire856 <<< wire856)))));
  assign wire860 = {wire841, wire844};
  assign wire861 = ((-(~|$unsigned((reg853 >> reg849)))) ?
                       ((reg849[(5'h13):(1'h1)] <<< wire857[(1'h0):(1'h0)]) & $signed($signed(reg850))) : $unsigned((^(wire842 ?
                           $unsigned(wire858) : $unsigned(reg855)))));
  assign wire862 = ({($signed(reg849[(5'h12):(3'h7)]) == $unsigned((wire860 ?
                               reg848 : reg848))),
                           (reg851 && (7'h4b))} ?
                       (~|wire861) : (^~reg847[(1'h0):(1'h0)]));
  assign wire863 = (($signed((~^(wire861 ?
                           wire845 : (8'h9e)))) >> ($signed((~|wire839)) ?
                           $signed(((8'hb6) ?
                               wire842 : (8'ha3))) : $signed($signed((7'h4e))))) ?
                       ({wire844,
                           ((~|wire842) ~^ (wire862 ~^ reg851))} && {wire842[(5'h10):(3'h6)]}) : ((~&wire844) <= $signed($signed({wire839}))));
  assign wire864 = (~$signed(((+wire841) ?
                       (+$unsigned(reg848)) : (((8'hb6) ? wire854 : wire839) ?
                           {wire862} : (7'h44)))));
  always
    @(posedge clk) begin
      if (({$signed({wire857, $signed(reg846)}),
          {(reg855[(3'h6):(2'h3)] != (~&wire843)),
              $unsigned($unsigned(reg851))}} ~^ $signed(wire859[(3'h5):(2'h2)])))
        begin
          if (($unsigned(wire856[(5'h11):(5'h10)]) ?
              {$unsigned($unsigned((reg852 & wire842)))} : ($unsigned($signed((!reg853))) ~^ wire858)))
            begin
              reg865 <= (reg851[(4'hb):(4'ha)] < ($signed(({reg852,
                  (8'hb9)} != $signed((7'h46)))) == (wire857 ?
                  ({(8'hbc)} ~^ $signed(wire840)) : {$signed(wire842)})));
            end
          else
            begin
              reg865 <= (wire859[(4'h8):(3'h5)] << ($unsigned((reg855 ?
                  (-wire863) : reg846)) + (($signed(wire839) >>> (~&(8'ha4))) ^ $unsigned({reg853}))));
              reg866 <= (~|$unsigned(((~{(8'hab), wire842}) ?
                  reg865 : wire840)));
              reg867 <= (~|(((wire863[(4'ha):(2'h3)] ?
                          $unsigned((8'hb8)) : reg849) ?
                      reg847 : (-$signed(wire860))) ?
                  (8'h9f) : (~&(^~reg865))));
              reg868 <= (8'ha5);
              reg869 <= ($signed(wire840[(3'h6):(3'h5)]) | reg853);
            end
          if ((8'ha9))
            begin
              reg870 <= $unsigned((+wire861[(4'hc):(3'h4)]));
              reg871 <= {$signed((!$signed(wire844)))};
              reg872 <= $unsigned({wire856, wire845[(3'h6):(3'h5)]});
            end
          else
            begin
              reg870 <= wire864[(3'h7):(3'h7)];
              reg871 <= reg850;
              reg872 <= ($unsigned((~^$signed($unsigned(reg846)))) ?
                  (~^$signed(wire857)) : ($signed($signed((~&wire857))) ?
                      reg846[(2'h2):(2'h2)] : ($signed({reg855, wire860}) ?
                          $unsigned(reg851) : (+$signed(wire861)))));
              reg873 <= reg852;
            end
          if (wire854)
            begin
              reg874 <= (reg868[(3'h7):(3'h5)] << (reg849 + (((~^reg855) <<< $unsigned(reg847)) != reg847[(2'h3):(1'h1)])));
              reg875 <= (wire844[(2'h3):(1'h0)] ?
                  wire859[(3'h5):(1'h1)] : $unsigned(({(~&wire859)} == $unsigned($signed(reg873)))));
              reg876 <= $unsigned($unsigned((^wire862[(5'h13):(3'h7)])));
              reg877 <= {(+(~&wire843)), (~reg876[(5'h11):(3'h6)])};
              reg878 <= (-reg851[(5'h1a):(3'h6)]);
            end
          else
            begin
              reg874 <= (wire845 ? wire861 : wire856);
              reg875 <= ({{((wire840 * (7'h40)) ~^ (8'ha4))}} <= $unsigned(wire862[(1'h0):(1'h0)]));
              reg876 <= $signed($unsigned({{(|reg872)}}));
              reg877 <= (8'ha5);
              reg878 <= (((~&$signed({reg866})) ?
                  (($unsigned(reg868) & $unsigned(wire861)) ?
                      reg850[(1'h0):(1'h0)] : reg850) : $signed((^$signed((7'h4e))))) * $signed(reg869[(1'h1):(1'h0)]));
            end
          if (reg874[(5'h11):(4'h8)])
            begin
              reg879 <= ((|(^reg865[(5'h1a):(4'ha)])) || ((wire844[(1'h1):(1'h1)] & $signed(wire859)) ~^ ($unsigned($signed(wire844)) | wire861[(4'hc):(4'h8)])));
              reg880 <= (-$unsigned($signed((~&(+reg851)))));
              reg881 <= {(wire863[(2'h3):(1'h0)] <= ($signed(wire863[(4'ha):(4'ha)]) + {(reg869 ^~ reg867)})),
                  reg869};
              reg882 <= wire856;
            end
          else
            begin
              reg879 <= reg881;
              reg880 <= reg869[(3'h5):(2'h3)];
              reg881 <= $signed(reg850[(5'h13):(4'hf)]);
              reg882 <= $signed((((-(^wire860)) ?
                  $signed((reg868 ^~ reg879)) : (~^$unsigned((7'h42)))) + (-{((8'had) < reg874),
                  (~&(8'hab))})));
              reg883 <= reg866[(4'h8):(3'h5)];
            end
        end
      else
        begin
          reg865 <= reg879;
        end
      reg884 <= reg850;
      if ($unsigned(((8'ha7) ?
          $signed((7'h4b)) : {{(wire842 >= wire845), wire859[(2'h3):(2'h3)]}})))
        begin
          if (wire861)
            begin
              reg885 <= $unsigned((reg868[(4'h8):(3'h5)] ?
                  (((wire859 * reg852) + (7'h41)) != {reg870[(5'h12):(4'h8)]}) : reg872));
              reg886 <= (reg851[(1'h1):(1'h0)] ?
                  {wire845,
                      {wire857,
                          reg875[(2'h2):(1'h0)]}} : ((-(&$unsigned((8'ha6)))) | $unsigned({(^~reg865)})));
            end
          else
            begin
              reg885 <= {{({(reg874 * reg885)} ^ $unsigned($unsigned(wire860))),
                      wire842},
                  (({(^(8'hb9))} && $signed($signed(reg867))) << wire854)};
              reg886 <= (&$unsigned({reg881, $unsigned($unsigned((7'h4d)))}));
            end
          reg887 <= (~|wire845);
          reg888 <= {reg866[(2'h2):(1'h1)], wire860};
        end
      else
        begin
          if ({reg846, {reg868}})
            begin
              reg885 <= ((|($signed({reg885}) >= (reg871[(2'h2):(1'h0)] ?
                  (wire842 ? reg881 : reg870) : (reg873 ?
                      (8'hb3) : reg867)))) == ((($signed(reg868) ?
                      (^wire840) : (wire860 ?
                          reg883 : wire863)) << $signed((reg880 && reg846))) ?
                  (((reg881 < wire864) ?
                      reg869[(2'h2):(1'h1)] : (|reg870)) | $unsigned(reg867[(3'h5):(3'h5)])) : (~|{(|(8'hb5))})));
              reg886 <= (~{$unsigned(reg873)});
              reg887 <= reg877[(3'h5):(3'h4)];
            end
          else
            begin
              reg885 <= $signed(reg855);
              reg886 <= wire842[(5'h19):(5'h13)];
            end
          if (reg871[(2'h2):(1'h0)])
            begin
              reg888 <= $signed({(~&($unsigned(reg886) >>> wire861[(1'h1):(1'h1)])),
                  $signed($signed((~|reg883)))});
              reg889 <= $signed($signed(((wire844 >> $signed(reg875)) ?
                  (reg876 | {wire859}) : (wire845[(2'h3):(1'h1)] ?
                      (~|(7'h44)) : reg874))));
            end
          else
            begin
              reg888 <= (+wire859);
              reg889 <= $unsigned((reg882[(4'hc):(3'h4)] << ($signed((reg888 ?
                  reg885 : reg874)) == ((8'ha6) ? reg884 : {reg885, reg850}))));
              reg890 <= (~&reg885);
              reg891 <= reg847;
              reg892 <= ($unsigned(((reg886 >> (reg872 ? reg846 : (7'h41))) ?
                      (~wire863) : $unsigned((8'hbc)))) ?
                  reg890 : reg891);
              reg893 <= {((reg874 > reg848[(2'h2):(2'h2)]) ^ ($unsigned(((8'ha9) ?
                          wire839 : reg889)) ?
                      (((8'ha0) ?
                          (8'ha7) : reg868) << reg889[(4'hf):(4'he)]) : wire843)),
                  ((reg888[(1'h0):(1'h0)] << reg875[(1'h0):(1'h0)]) ?
                      $unsigned((reg872 ?
                          $unsigned(reg886) : wire841[(3'h7):(1'h0)])) : reg885[(2'h2):(2'h2)])};
            end
          if ((!$unsigned(wire862)))
            begin
              reg894 <= (reg892 ?
                  reg847 : {(($signed(reg873) + (~reg884)) ?
                          (wire843 || reg852) : reg870[(3'h7):(1'h0)]),
                      ({$unsigned(wire840), $unsigned(reg855)} ?
                          ({reg886,
                              wire842} || $signed(reg890)) : (wire864[(3'h4):(2'h3)] ?
                              reg891[(5'h12):(4'he)] : $signed(reg848)))});
              reg895 <= reg870;
              reg896 <= $signed(reg846[(3'h5):(1'h0)]);
              reg897 <= {reg886[(3'h7):(3'h7)]};
              reg898 <= ((^~(reg866 ?
                  $unsigned({reg868}) : $unsigned($unsigned(reg897)))) == wire862);
              reg899 <= $unsigned(reg881);
            end
          else
            begin
              reg894 <= ($signed(((wire845 || $signed(wire841)) << ($unsigned(reg872) ?
                      reg877 : wire862[(3'h6):(3'h5)]))) ?
                  ((^($unsigned(wire844) ~^ $signed(wire841))) >> ($signed(reg871) << wire845)) : ($unsigned($signed((-wire844))) ?
                      reg847[(1'h1):(1'h0)] : (($signed(reg886) ?
                          $signed((8'ha5)) : (reg876 ?
                              reg897 : wire840)) ^~ $unsigned((~^reg898)))));
              reg895 <= reg891[(3'h6):(1'h1)];
              reg896 <= (reg884[(5'h16):(4'hb)] ^ reg873);
              reg897 <= $unsigned(wire845);
              reg898 <= (!(reg897 == reg891[(5'h11):(4'h8)]));
              reg899 <= reg866;
            end
          if ((reg872[(5'h14):(1'h1)] != $signed($unsigned(reg883[(2'h2):(1'h0)]))))
            begin
              reg900 <= ((reg885 ?
                  $unsigned(reg897) : {(~^reg883[(4'hc):(3'h6)]),
                      ($signed(reg896) <<< $signed(reg873))}) >> wire859);
              reg901 <= $signed(wire858);
            end
          else
            begin
              reg900 <= (8'hb9);
              reg901 <= (((8'ha6) ?
                      ({(reg883 ?
                              wire844 : reg894)} - $unsigned(wire859)) : (($signed(reg897) <= reg885[(3'h4):(2'h3)]) ?
                          $signed((~&reg882)) : reg900)) ?
                  {$unsigned(($unsigned((7'h40)) ?
                          $unsigned(reg900) : (8'ha3)))} : (-(~|reg874[(4'ha):(3'h5)])));
              reg902 <= (+$unsigned($signed(((reg847 || reg851) ?
                  $signed(reg897) : wire862))));
              reg903 <= {reg898, (|(~&({wire857} && (~&reg850))))};
            end
          if ((+$unsigned(reg866)))
            begin
              reg904 <= reg855[(1'h0):(1'h0)];
              reg905 <= {(~|(^(reg876[(4'h8):(3'h5)] ?
                      (reg897 ? reg855 : (8'hac)) : (reg855 == reg848))))};
            end
          else
            begin
              reg904 <= $unsigned((^~wire858[(4'hb):(3'h4)]));
              reg905 <= (reg901 ?
                  ($signed(((^~reg851) ?
                      (^~reg866) : wire839[(4'ha):(2'h2)])) ~^ (8'ha5)) : $unsigned((reg852[(2'h3):(2'h2)] | reg887[(4'h9):(2'h2)])));
            end
        end
    end
  assign wire906 = wire841;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module689  (y, clk, wire694, wire693, wire692, wire691, wire690);
  output wire [(32'h75c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire694;
  input wire signed [(4'hf):(1'h0)] wire693;
  input wire [(5'h19):(1'h0)] wire692;
  input wire signed [(3'h5):(1'h0)] wire691;
  input wire signed [(2'h2):(1'h0)] wire690;
  wire signed [(4'hd):(1'h0)] wire832;
  wire [(5'h11):(1'h0)] wire831;
  wire [(5'h14):(1'h0)] wire830;
  wire signed [(5'h18):(1'h0)] wire829;
  wire [(2'h2):(1'h0)] wire778;
  wire [(5'h15):(1'h0)] wire777;
  wire signed [(2'h3):(1'h0)] wire776;
  wire signed [(3'h6):(1'h0)] wire775;
  wire signed [(3'h4):(1'h0)] wire774;
  wire signed [(5'h17):(1'h0)] wire768;
  wire signed [(5'h1a):(1'h0)] wire767;
  wire [(2'h2):(1'h0)] wire766;
  wire signed [(5'h14):(1'h0)] wire765;
  wire signed [(5'h15):(1'h0)] wire762;
  wire signed [(3'h7):(1'h0)] wire761;
  wire [(4'hb):(1'h0)] wire760;
  wire signed [(3'h6):(1'h0)] wire759;
  wire signed [(5'h13):(1'h0)] wire758;
  wire [(3'h5):(1'h0)] wire757;
  reg signed [(3'h5):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg826 = (1'h0);
  reg [(3'h7):(1'h0)] reg825 = (1'h0);
  reg [(2'h2):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg823 = (1'h0);
  reg [(4'he):(1'h0)] reg822 = (1'h0);
  reg [(3'h4):(1'h0)] reg821 = (1'h0);
  reg [(5'h11):(1'h0)] reg820 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg818 = (1'h0);
  reg [(5'h12):(1'h0)] reg817 = (1'h0);
  reg [(5'h14):(1'h0)] reg816 = (1'h0);
  reg [(5'h18):(1'h0)] reg815 = (1'h0);
  reg [(3'h7):(1'h0)] reg814 = (1'h0);
  reg [(2'h2):(1'h0)] reg813 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg811 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg810 = (1'h0);
  reg [(5'h18):(1'h0)] reg809 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg808 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg807 = (1'h0);
  reg [(5'h18):(1'h0)] reg806 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg805 = (1'h0);
  reg [(3'h7):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg803 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg802 = (1'h0);
  reg [(4'h8):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg800 = (1'h0);
  reg [(5'h12):(1'h0)] reg799 = (1'h0);
  reg [(4'ha):(1'h0)] reg798 = (1'h0);
  reg [(5'h15):(1'h0)] reg797 = (1'h0);
  reg [(5'h12):(1'h0)] reg796 = (1'h0);
  reg [(3'h4):(1'h0)] reg795 = (1'h0);
  reg [(5'h1a):(1'h0)] reg794 = (1'h0);
  reg signed [(4'he):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg791 = (1'h0);
  reg [(3'h5):(1'h0)] reg790 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg789 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg788 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg787 = (1'h0);
  reg [(5'h13):(1'h0)] reg786 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg785 = (1'h0);
  reg [(4'h8):(1'h0)] reg784 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg783 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg782 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg780 = (1'h0);
  reg [(4'hb):(1'h0)] reg779 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg773 = (1'h0);
  reg [(4'hd):(1'h0)] reg772 = (1'h0);
  reg [(5'h11):(1'h0)] reg771 = (1'h0);
  reg [(5'h14):(1'h0)] reg770 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg769 = (1'h0);
  reg [(2'h2):(1'h0)] reg764 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg763 = (1'h0);
  reg [(5'h12):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg755 = (1'h0);
  reg [(4'h8):(1'h0)] reg754 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg753 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg752 = (1'h0);
  reg [(4'ha):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg750 = (1'h0);
  reg [(4'hb):(1'h0)] reg749 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg748 = (1'h0);
  reg [(5'h10):(1'h0)] reg747 = (1'h0);
  reg [(2'h3):(1'h0)] reg746 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg745 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg744 = (1'h0);
  reg [(5'h10):(1'h0)] reg743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg742 = (1'h0);
  reg [(3'h7):(1'h0)] reg741 = (1'h0);
  reg [(4'h9):(1'h0)] reg740 = (1'h0);
  reg [(3'h4):(1'h0)] reg739 = (1'h0);
  reg [(3'h6):(1'h0)] reg738 = (1'h0);
  reg [(2'h2):(1'h0)] reg737 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg736 = (1'h0);
  reg [(4'h9):(1'h0)] reg735 = (1'h0);
  reg [(5'h18):(1'h0)] reg734 = (1'h0);
  reg [(5'h12):(1'h0)] reg733 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg732 = (1'h0);
  reg [(3'h5):(1'h0)] reg731 = (1'h0);
  reg [(3'h4):(1'h0)] reg730 = (1'h0);
  reg [(5'h18):(1'h0)] reg729 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg727 = (1'h0);
  reg [(4'hb):(1'h0)] reg726 = (1'h0);
  reg [(5'h14):(1'h0)] reg725 = (1'h0);
  reg [(4'hf):(1'h0)] reg724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg723 = (1'h0);
  reg [(5'h14):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg721 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg720 = (1'h0);
  reg [(5'h10):(1'h0)] reg719 = (1'h0);
  reg [(4'hf):(1'h0)] reg718 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg717 = (1'h0);
  reg [(4'ha):(1'h0)] reg716 = (1'h0);
  reg [(2'h2):(1'h0)] reg715 = (1'h0);
  reg [(2'h2):(1'h0)] reg714 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg713 = (1'h0);
  reg [(3'h4):(1'h0)] reg712 = (1'h0);
  reg [(5'h1a):(1'h0)] reg711 = (1'h0);
  reg [(5'h17):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg709 = (1'h0);
  reg [(5'h11):(1'h0)] reg708 = (1'h0);
  reg [(2'h3):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg706 = (1'h0);
  reg [(4'ha):(1'h0)] reg705 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg704 = (1'h0);
  reg [(5'h17):(1'h0)] reg703 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg702 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg701 = (1'h0);
  reg [(5'h12):(1'h0)] reg700 = (1'h0);
  reg [(5'h14):(1'h0)] reg699 = (1'h0);
  reg [(5'h13):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg697 = (1'h0);
  reg [(5'h18):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg695 = (1'h0);
  assign y = {wire832,
                 wire831,
                 wire830,
                 wire829,
                 wire778,
                 wire777,
                 wire776,
                 wire775,
                 wire774,
                 wire768,
                 wire767,
                 wire766,
                 wire765,
                 wire762,
                 wire761,
                 wire760,
                 wire759,
                 wire758,
                 wire757,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg769,
                 reg764,
                 reg763,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 reg695,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((&wire693[(2'h3):(2'h3)]))
        begin
          if ($signed((wire692[(2'h3):(1'h0)] > wire694)))
            begin
              reg695 <= wire692;
              reg696 <= ((8'hac) + (($unsigned((wire693 < wire693)) | $unsigned((^(8'hb4)))) == (($signed((8'ha5)) ?
                      wire690 : reg695) ?
                  (|{(8'hbf), reg695}) : (~&$unsigned(wire691)))));
              reg697 <= reg696;
            end
          else
            begin
              reg695 <= $signed($unsigned(($signed($unsigned(reg695)) == $unsigned($signed(wire692)))));
              reg696 <= reg697;
              reg697 <= $unsigned(wire690[(1'h0):(1'h0)]);
              reg698 <= ($signed(wire693[(4'ha):(2'h3)]) >>> wire691[(3'h4):(2'h2)]);
              reg699 <= reg695;
              reg700 <= (reg697 ?
                  wire692[(2'h3):(2'h2)] : ((~|(~$unsigned(wire692))) + reg696[(5'h12):(1'h0)]));
            end
          reg701 <= (7'h4a);
          if ((+$signed(((~$signed(wire692)) ?
              reg700[(2'h2):(1'h0)] : $unsigned((~wire691))))))
            begin
              reg702 <= ((|$signed($unsigned((-reg696)))) ?
                  {$unsigned($unsigned($unsigned(wire692))),
                      reg699} : $signed((reg695[(1'h0):(1'h0)] ^~ reg695)));
              reg703 <= reg699;
              reg704 <= ((reg700 >>> $signed((~&reg702))) ?
                  $signed((-{reg698,
                      {(8'hb7), reg702}})) : $unsigned(reg700[(2'h2):(1'h1)]));
              reg705 <= $signed((8'hb4));
            end
          else
            begin
              reg702 <= ((reg697[(3'h4):(3'h4)] != $signed(reg697)) ?
                  $signed($unsigned(reg698[(3'h4):(1'h0)])) : $signed($signed(({wire692,
                      wire691} > (~|reg701)))));
              reg703 <= $signed(wire693[(2'h3):(2'h2)]);
              reg704 <= reg698[(3'h7):(3'h6)];
              reg705 <= (|({(^~(~&reg704)), (reg696 == reg702)} ?
                  ($signed($signed(reg700)) ?
                      {(wire690 >> wire691)} : (|$signed((8'ha0)))) : $unsigned(($unsigned(reg696) ~^ $signed(wire690)))));
              reg706 <= wire692;
              reg707 <= {(($signed($unsigned((8'h9c))) << ((wire694 ^~ reg696) ?
                          {reg697} : $unsigned((8'hb0)))) ?
                      (reg704[(1'h0):(1'h0)] & $signed(wire692[(2'h2):(1'h0)])) : wire694)};
            end
          reg708 <= (~|$unsigned($unsigned(reg695[(4'h8):(2'h2)])));
        end
      else
        begin
          if ((reg696 << (^~reg702)))
            begin
              reg695 <= $signed($signed(reg699));
            end
          else
            begin
              reg695 <= (!$unsigned((($signed((8'hab)) <<< wire692) ?
                  wire694[(3'h6):(3'h5)] : $unsigned((|(8'hb4))))));
            end
          if (($unsigned((((~reg703) + (reg696 ? (8'hb3) : reg703)) ?
              (~&(reg707 ?
                  (7'h41) : reg705)) : reg699)) >>> $signed((wire690 * ((reg698 ^~ wire693) ?
              $signed(reg707) : (reg705 ? wire694 : wire693))))))
            begin
              reg696 <= $signed($signed(wire690[(2'h2):(1'h1)]));
            end
          else
            begin
              reg696 <= $signed(($unsigned(wire693[(4'he):(3'h5)]) ?
                  reg698[(4'hc):(3'h5)] : (reg696[(5'h11):(4'h9)] >>> $unsigned(reg701))));
              reg697 <= (((reg695 != $signed($signed(reg698))) == wire690[(1'h0):(1'h0)]) ?
                  ($signed(reg703) && ((|reg700[(4'hf):(3'h6)]) && $unsigned((reg706 ?
                      reg696 : wire694)))) : (~^((+$signed(reg698)) || $signed((reg695 ?
                      reg708 : reg705)))));
              reg698 <= $signed(((reg701[(3'h6):(3'h6)] + (((8'hb9) ?
                      wire690 : (8'ha8)) * wire690[(1'h1):(1'h1)])) ?
                  $unsigned(reg706) : (wire690 ?
                      {{reg708}} : $unsigned((|wire690)))));
              reg699 <= reg702;
              reg700 <= (+{$unsigned($signed((reg695 ? reg703 : reg706))),
                  ((8'ha6) ~^ ((reg698 != reg704) ^~ $unsigned(wire691)))});
              reg701 <= ($unsigned($signed(wire694[(1'h0):(1'h0)])) != $signed(($signed((wire693 ?
                      reg704 : reg698)) ?
                  (+(~reg696)) : ($unsigned(wire690) << {reg705}))));
            end
          reg702 <= wire691;
        end
      if (reg697[(4'h8):(3'h4)])
        begin
          if (((~|((wire693 >>> wire692) ?
                  ((~&reg698) ? $unsigned(wire693) : wire694) : reg708)) ?
              reg698 : $unsigned($unsigned(reg708[(4'hf):(4'hd)]))))
            begin
              reg709 <= reg701[(3'h4):(1'h1)];
              reg710 <= {$unsigned($unsigned((~^$signed(reg701))))};
            end
          else
            begin
              reg709 <= $signed((8'hbb));
            end
        end
      else
        begin
          if ((reg703 << $unsigned((!(reg701[(2'h2):(1'h0)] ?
              ((8'ha5) << reg695) : (~|reg707))))))
            begin
              reg709 <= {{reg700[(5'h12):(4'hb)],
                      {((wire691 == (8'hab)) ?
                              $signed((7'h49)) : $unsigned(reg709)),
                          $signed((wire691 ? reg701 : wire693))}},
                  ((reg700 ?
                          ((~reg703) >>> (~reg706)) : $unsigned($unsigned(reg705))) ?
                      ($signed(reg695[(4'he):(1'h1)]) | wire694[(1'h0):(1'h0)]) : $signed($signed($unsigned((8'hb4)))))};
              reg710 <= (+reg699[(4'hb):(2'h3)]);
              reg711 <= ($signed(reg707[(2'h3):(2'h2)]) << ($signed(reg699) ?
                  {((+(8'hb6)) ? $unsigned(reg695) : $unsigned(reg708)),
                      reg707} : {(~^{reg701, reg704})}));
            end
          else
            begin
              reg709 <= $unsigned($unsigned((8'hb3)));
              reg710 <= $unsigned(reg698);
              reg711 <= reg710[(5'h17):(5'h12)];
              reg712 <= ($signed((reg702 ?
                  $unsigned($signed(reg709)) : $signed((!wire690)))) ^ $unsigned(reg699[(2'h2):(1'h0)]));
              reg713 <= ((^~$unsigned(((~^reg701) ?
                  (wire694 ?
                      reg712 : (8'hbb)) : (8'ha9)))) >>> (~|(&(wire694 || reg699))));
            end
          if ($signed((~^($signed((8'hab)) ?
              ((reg705 ? wire693 : wire690) ^ (reg698 ?
                  reg702 : reg712)) : $signed(wire692)))))
            begin
              reg714 <= (^(((8'hbc) || reg697[(4'hf):(3'h7)]) ?
                  reg710[(4'he):(3'h7)] : reg697));
              reg715 <= $signed(({$signed($signed(reg706)),
                      reg696[(4'he):(3'h4)]} ?
                  $signed($unsigned(reg698)) : reg702));
              reg716 <= (8'ha0);
              reg717 <= $unsigned((~|$unsigned(reg716[(3'h6):(2'h3)])));
              reg718 <= reg716;
            end
          else
            begin
              reg714 <= ((reg701 < (reg704[(1'h1):(1'h1)] + wire693)) == reg698[(4'hc):(3'h6)]);
              reg715 <= (7'h4d);
              reg716 <= $unsigned($unsigned($signed(reg695[(1'h0):(1'h0)])));
              reg717 <= ((8'hb8) ? reg715 : reg700[(1'h0):(1'h0)]);
              reg718 <= {$signed(reg716), (|reg711)};
            end
          reg719 <= $unsigned($unsigned((^~reg699)));
          reg720 <= {$signed(reg704)};
          if ({$unsigned((^(!{reg698, reg703})))})
            begin
              reg721 <= (reg698 ?
                  (($signed((wire691 && wire692)) ?
                      $signed({reg720}) : (~(reg716 >>> (8'h9f)))) == {{(wire693 ?
                              reg720 : wire692)}}) : $unsigned($unsigned(((wire693 == reg708) == (-reg714)))));
              reg722 <= (reg707[(1'h1):(1'h0)] ?
                  reg716[(2'h2):(2'h2)] : reg698);
              reg723 <= ((~|((8'hb5) * $signed(reg718[(4'h9):(4'h8)]))) ?
                  ($unsigned((~&$signed(reg711))) ^~ $unsigned(wire693)) : {(^$unsigned((~&wire693)))});
              reg724 <= $unsigned($signed(reg719[(4'ha):(3'h6)]));
              reg725 <= (reg696 ?
                  $unsigned($signed((reg708 <<< $signed(reg704)))) : ($unsigned(reg715) + ((&(+reg721)) ?
                      $unsigned($signed(reg719)) : ((reg708 != reg702) ?
                          ((8'ha3) ? reg717 : reg698) : reg714))));
            end
          else
            begin
              reg721 <= ({$signed($signed($unsigned(reg698)))} ?
                  reg707 : $signed($unsigned($signed((reg702 >>> reg697)))));
              reg722 <= ($unsigned(((reg709 - {reg702,
                  (8'h9e)}) <<< ($unsigned(reg700) < (|reg708)))) & {reg718[(3'h5):(2'h3)]});
              reg723 <= {reg722, reg715[(1'h0):(1'h0)]};
              reg724 <= reg719[(3'h5):(1'h0)];
              reg725 <= reg700[(5'h10):(2'h3)];
              reg726 <= reg711[(5'h16):(3'h5)];
            end
          reg727 <= reg711;
        end
      if (reg705)
        begin
          if ({$unsigned(($signed(reg696) == $signed(reg722)))})
            begin
              reg728 <= $signed(((!(-((7'h43) ? reg709 : wire694))) ?
                  (reg716[(3'h7):(1'h0)] ?
                      (reg695 ?
                          (reg698 ?
                              (7'h4d) : (8'hb0)) : reg710) : reg727[(4'h8):(3'h6)]) : $unsigned((^reg727))));
              reg729 <= (~&$signed((({reg697} ? $signed((7'h42)) : (~|reg726)) ?
                  (reg695[(4'hd):(4'h9)] ?
                      wire690[(2'h2):(1'h0)] : $signed(wire694)) : $unsigned($unsigned(reg707)))));
              reg730 <= ((^reg703) ~^ $signed($unsigned($unsigned(reg722[(3'h6):(3'h4)]))));
              reg731 <= (~^((^~$signed({reg712})) << reg712[(2'h2):(1'h1)]));
              reg732 <= reg699[(4'h9):(3'h7)];
              reg733 <= $unsigned($unsigned(reg724[(2'h3):(1'h0)]));
            end
          else
            begin
              reg728 <= ((!$signed($unsigned($unsigned(reg730)))) | reg727);
              reg729 <= $unsigned((($signed($signed(wire694)) + $signed((-reg715))) > $unsigned((7'h41))));
              reg730 <= ((8'hbd) ? $unsigned($signed(reg733)) : (8'hb0));
              reg731 <= reg727;
              reg732 <= {$unsigned((reg721 ?
                      ((reg715 ? wire692 : reg699) ?
                          (-wire690) : (~reg711)) : (^$unsigned(reg702)))),
                  (($unsigned((8'hb4)) ?
                      $unsigned(wire690) : $signed((reg728 >= (8'ha8)))) ^~ reg730)};
            end
        end
      else
        begin
          if ($signed(wire690))
            begin
              reg728 <= $signed($unsigned((reg716 ?
                  reg714[(1'h1):(1'h1)] : {$signed((8'h9f)), (-reg728)})));
              reg729 <= (~^(&{wire693}));
              reg730 <= ((8'hb8) ? reg695 : reg725[(4'hf):(2'h3)]);
              reg731 <= ({reg711[(2'h3):(1'h1)]} ?
                  reg717[(1'h0):(1'h0)] : (reg726 << (^((reg704 >> reg721) ?
                      (reg700 << reg728) : (~|wire694)))));
              reg732 <= ((+((7'h48) + reg732[(3'h4):(2'h3)])) || ((~|reg733[(2'h3):(1'h1)]) < ({reg719[(3'h4):(1'h1)]} ?
                  $unsigned($unsigned(reg706)) : reg719[(4'hc):(4'h9)])));
            end
          else
            begin
              reg728 <= reg717[(4'he):(4'hd)];
            end
          if ((~reg708))
            begin
              reg733 <= $unsigned({$signed($signed(reg705[(1'h0):(1'h0)])),
                  ($signed((wire694 >> reg711)) ?
                      reg723 : ((reg733 | wire690) ?
                          (reg716 ? (7'h4b) : (8'hb2)) : $unsigned(reg720)))});
              reg734 <= (($unsigned(((wire694 ^ (8'hba)) >= (|reg730))) >= (~(reg709[(2'h3):(2'h2)] ?
                  reg719 : $signed(reg722)))) > $unsigned((|{reg711,
                  $unsigned(reg715)})));
            end
          else
            begin
              reg733 <= ((wire692[(4'hb):(3'h5)] ?
                      ((reg725[(5'h14):(5'h14)] >>> (!reg710)) ?
                          (!reg730[(3'h4):(2'h2)]) : {((8'hbd) >> reg701),
                              reg723[(1'h0):(1'h0)]}) : reg703) ?
                  {reg712} : ($unsigned(((~wire693) - $signed(wire691))) ?
                      $unsigned(((reg724 <= reg730) ~^ {reg713,
                          reg714})) : (({reg707} << $unsigned(reg703)) ?
                          {(|reg719)} : (~|$unsigned(reg733)))));
              reg734 <= reg708;
              reg735 <= ((!reg726) ?
                  ((reg715 * (reg714 ?
                      reg729[(1'h0):(1'h0)] : (reg733 >>> (8'hbd)))) & ($unsigned(wire692[(4'hb):(1'h0)]) ~^ ((reg717 ?
                      (7'h4e) : reg701) || (!reg723)))) : $signed(wire691));
              reg736 <= wire693[(4'ha):(4'h9)];
              reg737 <= (8'ha7);
              reg738 <= $signed($unsigned(((8'hba) ?
                  reg721[(5'h15):(1'h1)] : ((reg725 ?
                      reg724 : reg736) & (reg699 ? reg729 : reg717)))));
            end
          reg739 <= ($unsigned($signed({(reg704 | reg734)})) ?
              ((reg712 ? reg709[(4'he):(3'h6)] : (7'h4c)) ?
                  reg726 : ((~{reg735}) >> (&(~|reg717)))) : reg734);
          reg740 <= (~|reg727[(3'h6):(2'h3)]);
        end
      if (reg710[(4'h9):(3'h5)])
        begin
          reg741 <= (+$unsigned(reg708));
          if ((^{(8'hab), reg737[(1'h1):(1'h1)]}))
            begin
              reg742 <= reg703;
              reg743 <= $unsigned(reg739);
              reg744 <= reg739;
            end
          else
            begin
              reg742 <= {$signed($unsigned($unsigned($unsigned(reg713)))),
                  (($unsigned(reg732[(1'h1):(1'h0)]) ?
                          (&$signed(reg740)) : ((^reg743) * (|reg710))) ?
                      reg698[(3'h5):(2'h2)] : (+$unsigned($signed(reg714))))};
              reg743 <= (($signed(reg726[(4'h9):(4'h8)]) >= {{{reg711, reg714},
                          (wire692 ? reg698 : (7'h47))},
                      reg732[(1'h1):(1'h0)]}) ?
                  ((((reg744 && wire694) << {reg732}) - {$unsigned(reg734),
                          (reg741 ? reg714 : (8'hb2))}) ?
                      (reg697[(3'h5):(1'h1)] ?
                          {wire691[(3'h5):(3'h5)],
                              $signed(reg720)} : {reg742[(4'h9):(3'h5)]}) : reg730[(3'h4):(2'h2)]) : reg710[(2'h2):(1'h1)]);
              reg744 <= ((+reg725[(3'h7):(2'h2)]) ?
                  reg719[(4'hd):(4'ha)] : $signed(reg726));
              reg745 <= (~|(wire694 ?
                  (&$unsigned((reg698 <= reg702))) : reg695));
              reg746 <= ((reg698[(4'hf):(4'hd)] ?
                  (~$unsigned(reg704)) : $unsigned((+(|reg695)))) << {($unsigned(reg720) ?
                      $unsigned((reg734 >>> reg743)) : (+{(8'hac)})),
                  reg696[(5'h18):(5'h13)]});
            end
          if ($signed(({(~$signed((8'hbd)))} ?
              $signed({reg731[(2'h3):(1'h0)]}) : $signed(((~|reg703) ~^ $signed((8'hb6)))))))
            begin
              reg747 <= (7'h40);
              reg748 <= ({(~^(reg703 ?
                          {reg727} : ((8'h9d) ? reg722 : wire691))),
                      reg695[(2'h3):(2'h3)]} ?
                  (-$signed((-(-reg700)))) : reg734);
              reg749 <= (+$unsigned((|((-reg731) ? (-reg722) : {reg742}))));
              reg750 <= {$unsigned(reg724), reg721[(5'h11):(3'h6)]};
              reg751 <= $unsigned((|((reg743[(3'h5):(2'h3)] > (reg706 - reg750)) * $signed((reg723 ?
                  reg724 : reg739)))));
            end
          else
            begin
              reg747 <= (reg696[(2'h2):(1'h0)] ?
                  (~^reg741[(1'h0):(1'h0)]) : (((~(8'ha2)) ?
                      {$signed(reg718)} : (8'ha7)) && reg698));
              reg748 <= (reg744[(3'h7):(3'h6)] <<< reg728);
              reg749 <= $signed({($signed($signed((7'h4d))) ?
                      $signed((reg717 > (7'h47))) : ((+reg705) < (7'h41)))});
            end
          reg752 <= ((wire690 && reg723) > reg715);
          reg753 <= ((~(~&reg708)) == ($unsigned((~^(~|reg715))) ?
              {$signed(wire691)} : {(wire692[(1'h1):(1'h1)] ?
                      reg709 : reg738)}));
          reg754 <= (!(reg712[(2'h2):(1'h0)] >= reg726[(4'hb):(3'h7)]));
        end
      else
        begin
          reg741 <= ((+($signed($unsigned((8'ha1))) ?
                  $signed($unsigned((8'ha9))) : $unsigned(reg728[(4'hb):(4'h9)]))) ?
              reg739[(1'h0):(1'h0)] : {$signed(reg724[(1'h0):(1'h0)]),
                  $unsigned(wire690)});
          reg742 <= $unsigned(wire694[(3'h5):(1'h1)]);
          reg743 <= ($signed(reg702) ?
              reg724 : {$unsigned({reg716[(3'h4):(1'h0)],
                      reg737[(1'h0):(1'h0)]})});
          if ((reg723 ?
              $unsigned(reg731) : $signed(((~^reg705[(3'h5):(1'h1)]) ~^ ($signed(reg697) ^~ (7'h45))))))
            begin
              reg744 <= (wire691 >> reg701);
              reg745 <= ($signed((~|((-wire693) ? (~|reg750) : (~|reg730)))) ?
                  ((~&wire694[(2'h2):(2'h2)]) || reg703[(4'h8):(3'h6)]) : $unsigned(reg725[(5'h10):(4'he)]));
              reg746 <= ({(((reg702 ?
                          reg747 : reg726) == {(7'h4a)}) | $signed((reg730 ?
                          wire691 : wire691))),
                      ($signed($signed(reg727)) ?
                          reg751[(4'h8):(3'h4)] : $signed(((8'hb1) ?
                              (7'h42) : reg754)))} ?
                  (reg709[(3'h5):(2'h3)] ?
                      $signed($unsigned((reg720 >>> (7'h41)))) : $unsigned(reg702[(2'h3):(1'h0)])) : $signed($unsigned(((^reg700) + $signed((8'hb4))))));
            end
          else
            begin
              reg744 <= (~^reg730);
              reg745 <= (8'had);
              reg746 <= $unsigned(($unsigned(($unsigned(reg714) * reg697)) ^~ reg720[(4'h9):(3'h4)]));
              reg747 <= $unsigned((~&reg728));
              reg748 <= $signed((~&$signed(reg695)));
              reg749 <= reg730;
            end
          if (reg702)
            begin
              reg750 <= ((((~reg737) >= $signed(reg715)) | ($signed((reg730 >>> reg742)) == (+reg730[(1'h0):(1'h0)]))) ?
                  {$unsigned(($unsigned(reg724) != (|reg708)))} : $unsigned(reg698));
            end
          else
            begin
              reg750 <= $unsigned($signed((7'h42)));
              reg751 <= reg753;
              reg752 <= ($unsigned($unsigned($signed({reg733, reg705}))) ?
                  $unsigned($unsigned(reg747)) : reg752[(3'h6):(2'h3)]);
              reg753 <= (~&$unsigned(reg741[(1'h1):(1'h1)]));
              reg754 <= ($signed(wire694[(3'h7):(3'h6)]) >= (reg711[(5'h16):(3'h7)] == reg702[(2'h2):(1'h0)]));
              reg755 <= {{(~&((reg752 > reg754) - (wire691 ?
                          reg717 : reg703)))},
                  ($unsigned({reg722[(2'h3):(1'h1)],
                          (reg696 ? reg710 : reg707)}) ?
                      $signed($unsigned((reg716 ?
                          (8'ha1) : (7'h4c)))) : $signed($unsigned($signed((8'hbf)))))};
            end
          reg756 <= (+(((!$signed(reg725)) ?
              $unsigned(((8'ha6) >= reg707)) : ((reg749 ?
                  reg701 : reg731) ~^ {(7'h43)})) >>> reg748[(1'h0):(1'h0)]));
        end
    end
  assign wire757 = (($signed(reg696[(1'h0):(1'h0)]) ?
                       (reg722 << reg699) : (~|(-(reg708 ~^ reg713)))) <= reg712);
  assign wire758 = (^~reg720[(4'h9):(3'h5)]);
  assign wire759 = reg708;
  assign wire760 = $unsigned(reg737[(1'h1):(1'h1)]);
  assign wire761 = (|{(-((&reg730) <<< reg726)), {reg722}});
  assign wire762 = $signed($unsigned($signed(((reg714 ? wire694 : reg742) ?
                       $unsigned(reg707) : $signed((8'hb2))))));
  always
    @(posedge clk) begin
      reg763 <= ((((7'h4a) >> reg705) ?
              (reg754[(1'h1):(1'h0)] + (reg707[(1'h0):(1'h0)] || (wire758 <= wire762))) : (($signed(wire690) ?
                  (+wire757) : (reg706 ?
                      reg748 : (8'ha5))) ~^ $unsigned({reg704}))) ?
          wire691[(2'h2):(1'h0)] : (($unsigned((reg747 || reg751)) ?
                  reg725 : reg749[(4'ha):(4'h9)]) ?
              reg710 : reg742));
      reg764 <= reg747;
    end
  assign wire765 = ({(((reg740 ? wire693 : wire757) && reg729[(3'h4):(2'h3)]) ?
                               $signed($signed(reg723)) : ((reg721 >>> reg715) >= {reg730})),
                           reg708[(3'h5):(3'h5)]} ?
                       reg753[(3'h4):(2'h2)] : ({(8'h9f),
                           (!(^~reg718))} ^~ $signed({(reg719 ?
                               reg707 : (7'h47)),
                           (reg728 >= reg720)})));
  assign wire766 = (((!reg744[(3'h5):(3'h4)]) ~^ (((reg764 ?
                           reg709 : reg744) >= reg707) + ((~^reg718) ?
                           ((8'hb4) ? wire762 : (8'hb2)) : (-reg755)))) ?
                       (8'ha3) : (-(8'ha2)));
  assign wire767 = ($unsigned(reg701[(2'h3):(2'h2)]) ~^ (7'h44));
  assign wire768 = (^~{((!reg737[(2'h2):(2'h2)]) ?
                           wire765 : ($signed(wire767) > $signed((8'ha7))))});
  always
    @(posedge clk) begin
      if ((~^$signed(reg737[(1'h0):(1'h0)])))
        begin
          if (reg721)
            begin
              reg769 <= $unsigned($unsigned((wire761[(3'h5):(3'h4)] >> $signed((~^reg718)))));
              reg770 <= {reg732[(3'h4):(1'h1)],
                  (((&$unsigned((8'hba))) ?
                          ({reg748} >>> (reg739 ?
                              reg743 : reg708)) : ($unsigned(reg714) << (reg711 ?
                              wire767 : wire757))) ?
                      $unsigned(reg739) : ($signed((reg719 >>> reg755)) ^~ (^~reg703)))};
              reg771 <= $signed(({$signed(reg733[(3'h5):(1'h0)]),
                  reg714[(1'h0):(1'h0)]} == reg722));
              reg772 <= $unsigned($unsigned({{(-(7'h42))}}));
              reg773 <= wire762;
            end
          else
            begin
              reg769 <= (($signed(($signed(reg707) > (~reg699))) << reg716[(2'h3):(1'h0)]) * $signed(reg695[(1'h0):(1'h0)]));
              reg770 <= reg738[(2'h3):(1'h1)];
              reg771 <= (&$unsigned($signed(reg744)));
            end
        end
      else
        begin
          reg769 <= reg736;
          reg770 <= $unsigned((|((8'ha8) >> reg719)));
          reg771 <= (reg769 < ((((|wire759) ?
                  (^wire693) : $signed(reg710)) >>> (|(reg699 - wire757))) ?
              (({reg717, reg745} ?
                  (-reg704) : {wire692}) | reg725) : ($unsigned(reg703) ^~ $unsigned(reg703))));
        end
    end
  assign wire774 = ({(((-reg697) ? ((8'ha4) >= (8'hb6)) : reg732) < (7'h4a))} ?
                       (reg706[(3'h4):(2'h3)] <= reg745) : (|($signed((reg733 ?
                               wire765 : reg734)) ?
                           (^$signed(wire766)) : {wire692,
                               (reg704 ? reg716 : (7'h42))})));
  assign wire775 = {$unsigned(((~(~^reg726)) ?
                           ($unsigned((8'hb4)) | (wire774 ?
                               reg721 : wire761)) : wire768)),
                       ($unsigned($signed(reg729)) ?
                           ($unsigned($unsigned(reg701)) ?
                               ({reg746} << reg705[(4'ha):(4'ha)]) : reg744[(4'hb):(1'h0)]) : (+(reg763[(2'h3):(1'h0)] <= (-reg711))))};
  assign wire776 = $signed((^$unsigned(wire759)));
  assign wire777 = $signed(($unsigned(wire761) ?
                       reg707 : ((~|$signed(reg744)) ~^ $unsigned((reg706 + wire757)))));
  assign wire778 = (~&($signed(reg715[(1'h0):(1'h0)]) ?
                       (&(~&$signed(reg748))) : (reg763 ?
                           ((8'hb0) > $signed(reg712)) : $unsigned((reg725 ?
                               reg772 : reg742)))));
  always
    @(posedge clk) begin
      reg779 <= (7'h40);
      reg780 <= ((reg756[(4'hf):(3'h4)] >>> ((|(&reg745)) ?
          $unsigned($unsigned(wire767)) : ($signed(reg695) & reg769))) || $signed((^({reg722} >>> reg755))));
    end
  always
    @(posedge clk) begin
      reg781 <= reg698[(4'h8):(3'h6)];
      if (reg746)
        begin
          reg782 <= {(^(reg734 ?
                  $unsigned((reg780 ? reg704 : reg755)) : $signed((^~reg697)))),
              (8'ha2)};
          if (reg755[(5'h12):(5'h12)])
            begin
              reg783 <= $unsigned(reg723);
              reg784 <= reg720;
            end
          else
            begin
              reg783 <= reg732[(1'h0):(1'h0)];
            end
          if (((~^{$unsigned(reg716)}) && ($unsigned($signed($unsigned(reg714))) & $unsigned({(wire766 <= reg773),
              (7'h49)}))))
            begin
              reg785 <= $signed($signed((reg773[(4'hf):(3'h5)] ?
                  ($unsigned(wire692) ~^ (reg773 == reg717)) : reg716)));
              reg786 <= wire766[(1'h1):(1'h1)];
              reg787 <= ($signed($unsigned($unsigned((reg696 > reg706)))) ~^ reg730[(2'h2):(1'h0)]);
              reg788 <= ({(wire694 + ({reg782} <= (reg736 ? (8'h9f) : reg746))),
                  $unsigned($signed($signed(reg714)))} << $unsigned((^~reg716)));
              reg789 <= ((((^((7'h44) != reg772)) <<< ((^reg744) ?
                  reg780 : reg788[(4'ha):(1'h1)])) && $signed(($signed(reg770) - (reg755 != wire757)))) >= $unsigned($unsigned((|wire761))));
            end
          else
            begin
              reg785 <= ((((^~$signed((8'ha6))) >> reg769) ?
                  $signed($unsigned($unsigned(reg740))) : (&reg780[(2'h3):(2'h2)])) > ($unsigned((-reg720)) * (&(7'h4a))));
              reg786 <= ((wire768 ?
                  (~^$unsigned((wire767 << wire761))) : $signed($unsigned(reg744))) > wire693);
              reg787 <= (($unsigned(reg742[(4'hd):(3'h4)]) ?
                  {$signed(reg749),
                      (~|{reg752,
                          (8'hbd)})} : $signed((+reg738[(3'h5):(3'h5)]))) != {reg734});
              reg788 <= ((8'hbe) ?
                  reg703 : ((((~&reg700) * $unsigned(reg696)) ?
                          (~(^~(8'hb6))) : $unsigned((reg696 ?
                              reg714 : wire694))) ?
                      reg772[(3'h5):(3'h5)] : wire767[(5'h12):(4'h9)]));
              reg789 <= reg729;
            end
        end
      else
        begin
          if (wire767)
            begin
              reg782 <= reg704;
              reg783 <= ((((!wire690[(1'h1):(1'h0)]) - $signed((reg764 ?
                          (7'h4b) : reg733))) ?
                      $unsigned($signed($signed(reg769))) : {$unsigned(reg781[(2'h2):(1'h0)])}) ?
                  (($unsigned({reg740}) ?
                          reg763[(2'h2):(1'h1)] : reg784[(2'h2):(2'h2)]) ?
                      {reg719,
                          ($unsigned(wire759) || (^~reg752))} : ((8'hb4) << reg744[(5'h10):(4'hf)])) : wire691);
              reg784 <= reg783[(2'h2):(1'h0)];
              reg785 <= $signed({(($unsigned(reg749) ?
                      $signed((7'h44)) : $signed(reg695)) ^~ reg789[(4'hb):(3'h5)]),
                  (-((~^wire761) && reg736[(1'h0):(1'h0)]))});
            end
          else
            begin
              reg782 <= (^$unsigned(reg746[(1'h0):(1'h0)]));
              reg783 <= reg742[(1'h1):(1'h0)];
              reg784 <= $unsigned((~reg702));
              reg785 <= $signed(((reg731[(3'h5):(3'h4)] | ((7'h4d) < reg770[(2'h2):(1'h0)])) ?
                  {(|(reg745 << reg782)),
                      $unsigned((^reg784))} : {($signed(wire761) <= wire690[(2'h2):(1'h1)])}));
              reg786 <= $unsigned(wire760[(4'ha):(4'h8)]);
              reg787 <= $unsigned((|wire757));
            end
          if ({$signed(($signed(((8'h9d) <<< wire694)) ?
                  $unsigned((reg746 ? reg729 : reg697)) : ((reg696 >> (8'hac)) ?
                      $signed(reg749) : (reg717 + reg750))))})
            begin
              reg788 <= wire761[(3'h5):(1'h1)];
              reg789 <= ({(|reg741[(3'h4):(2'h2)])} << ($signed(($unsigned(reg748) ^ $unsigned(reg789))) ?
                  $unsigned($unsigned($unsigned(reg746))) : $unsigned(({reg780} && (8'ha4)))));
              reg790 <= reg737;
              reg791 <= $signed(reg698);
              reg792 <= $signed(reg725[(4'hf):(3'h7)]);
            end
          else
            begin
              reg788 <= ($unsigned(({$signed(reg704)} ?
                  ($unsigned(wire693) ?
                      (wire761 >> reg785) : reg717) : $signed(reg723))) ^~ wire768);
              reg789 <= reg730[(2'h2):(1'h1)];
            end
          reg793 <= (wire691 ?
              (wire766[(1'h1):(1'h0)] || ((-{reg727, reg745}) ?
                  $signed(reg745[(2'h3):(2'h3)]) : {reg717})) : wire761);
          if ($unsigned($unsigned({($signed(reg705) ?
                  ((8'ha0) * reg741) : (+reg783))})))
            begin
              reg794 <= (($unsigned(reg754) ?
                      $unsigned($unsigned(reg779[(3'h6):(3'h4)])) : (~^$signed({reg751}))) ?
                  (8'ha5) : ((7'h47) ?
                      reg779[(2'h2):(1'h0)] : (^(~$signed(reg730)))));
              reg795 <= ((~^{$signed(wire777[(4'hb):(2'h2)]),
                  reg790}) << ($unsigned($signed(reg734[(4'h9):(3'h6)])) ?
                  $unsigned($unsigned((wire774 ?
                      wire774 : reg712))) : ((8'hb0) ?
                      reg729 : $signed(reg735))));
              reg796 <= ($unsigned((((reg737 != (7'h4c)) ?
                      {reg793} : $unsigned(reg780)) ?
                  $unsigned((reg793 ?
                      reg724 : reg721)) : reg727[(5'h10):(3'h5)])) ^ reg782);
              reg797 <= $signed($unsigned(reg783[(1'h0):(1'h0)]));
            end
          else
            begin
              reg794 <= $unsigned(((!$signed(wire777)) ?
                  reg743 : $signed(reg702[(3'h5):(1'h1)])));
              reg795 <= $unsigned((~&(reg783[(3'h4):(3'h4)] ?
                  (reg706 ? (-reg743) : (reg744 >= reg709)) : {((8'ha8) ?
                          reg752 : (7'h4c)),
                      reg783[(2'h3):(1'h1)]})));
              reg796 <= (-$signed(reg739[(3'h4):(1'h0)]));
              reg797 <= (^(reg706[(5'h16):(3'h5)] ?
                  $signed((reg786[(5'h12):(5'h10)] && wire760[(3'h6):(2'h2)])) : $signed(wire691[(3'h5):(1'h0)])));
              reg798 <= (8'h9c);
              reg799 <= reg707;
            end
          reg800 <= $signed(reg724[(1'h1):(1'h0)]);
        end
      if ((&$unsigned(reg696)))
        begin
          if ((&$signed(wire774)))
            begin
              reg801 <= (+(((~&(&reg797)) ?
                  reg717[(1'h1):(1'h0)] : {{reg735, reg795},
                      reg718}) + {((8'hb9) ?
                      (reg745 ? (8'ha3) : reg782) : (reg796 ?
                          wire693 : reg726)),
                  wire774}));
              reg802 <= (reg715 ?
                  reg708[(3'h4):(2'h3)] : ((reg733[(3'h7):(2'h3)] | reg716) << reg792[(3'h4):(3'h4)]));
              reg803 <= reg726[(4'h8):(3'h4)];
              reg804 <= $unsigned(($signed((!reg752)) - $unsigned(reg787)));
              reg805 <= ((~^(wire692[(5'h17):(3'h5)] < $signed((^~reg751)))) ?
                  ((^~{$signed(reg718)}) + $unsigned(reg706[(4'hf):(2'h3)])) : (wire775 && reg748));
              reg806 <= (7'h4a);
            end
          else
            begin
              reg801 <= reg786[(4'he):(4'he)];
              reg802 <= wire762[(2'h2):(2'h2)];
            end
          if ((reg787[(1'h1):(1'h1)] << reg710))
            begin
              reg807 <= {$signed(wire778[(2'h2):(2'h2)])};
              reg808 <= ($signed((reg784 ?
                  ($signed(reg764) ?
                      $signed((7'h47)) : $signed(reg697)) : ($signed((8'hbf)) ?
                      {reg799, reg715} : (!reg709)))) > (reg795 ?
                  reg718[(2'h3):(2'h2)] : wire778[(1'h1):(1'h0)]));
            end
          else
            begin
              reg807 <= (reg796 ? reg748 : (&(8'ha7)));
              reg808 <= (~&$unsigned(reg735[(1'h0):(1'h0)]));
            end
          reg809 <= (!(~((&$signed((8'hbd))) ?
              $unsigned($signed(reg722)) : $unsigned(((8'ha4) <<< reg750)))));
        end
      else
        begin
          if ((~^$unsigned(wire774)))
            begin
              reg801 <= reg756;
              reg802 <= reg717[(5'h10):(4'h9)];
              reg803 <= (+(^~reg705[(4'h8):(1'h1)]));
              reg804 <= {reg734[(5'h18):(3'h6)], wire766};
            end
          else
            begin
              reg801 <= wire758[(4'hf):(4'h9)];
              reg802 <= ((~&$signed(((reg730 ?
                      wire768 : reg724) >= (~&reg802)))) ?
                  $unsigned(reg747[(5'h10):(2'h2)]) : $signed($unsigned(((reg781 <<< reg741) | reg785[(2'h3):(1'h0)]))));
              reg803 <= $signed((~((reg704[(5'h13):(4'hf)] <<< {reg710,
                  reg726}) + (reg807[(3'h6):(2'h2)] ?
                  (reg793 ^~ reg697) : $signed(wire777)))));
              reg804 <= ((reg755[(4'h8):(4'h8)] >>> $unsigned($signed((wire759 ?
                      (8'ha7) : reg708)))) ?
                  (^~(8'ha0)) : $unsigned((!$signed((reg695 ^ reg695)))));
              reg805 <= reg750;
              reg806 <= (~^reg702[(2'h2):(1'h1)]);
            end
          reg807 <= reg714[(1'h1):(1'h1)];
          if (((~|(~&reg726)) > $unsigned($signed((^reg705[(3'h4):(2'h2)])))))
            begin
              reg808 <= $signed($signed($unsigned($unsigned((reg785 ?
                  reg746 : wire778)))));
              reg809 <= ((wire692[(4'h9):(3'h5)] ?
                      $unsigned($unsigned($unsigned(wire777))) : (~&reg763[(3'h7):(3'h5)])) ?
                  {$signed((~&(reg742 ? reg771 : reg736))),
                      (reg800[(4'hb):(4'h8)] ~^ (^~$signed(reg729)))} : $unsigned($signed($signed($signed((8'ha9))))));
            end
          else
            begin
              reg808 <= reg771[(5'h11):(5'h11)];
              reg809 <= ({reg722[(2'h3):(2'h3)],
                  {(reg739 | wire762[(5'h13):(4'hc)]),
                      {$signed((7'h4d))}}} + ({$unsigned(reg773[(1'h0):(1'h0)]),
                  (((8'hb6) ? reg748 : reg745) ?
                      $signed(wire761) : reg721)} <<< (reg743 ?
                  (~reg738) : (~(~^reg700)))));
            end
          reg810 <= {(8'haf)};
          if (({((reg789 ? reg704 : (&reg726)) ?
                  $signed((reg763 ?
                      wire776 : reg730)) : wire777)} != reg710[(3'h7):(1'h0)]))
            begin
              reg811 <= $unsigned((!$unsigned(reg770[(4'hf):(4'hf)])));
              reg812 <= $unsigned({reg793});
              reg813 <= $signed(reg726);
              reg814 <= reg730;
              reg815 <= $signed((~&(~|(|reg795[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg811 <= (&reg805[(1'h0):(1'h0)]);
            end
        end
      if ((((-($unsigned(reg726) ? (7'h4e) : reg719)) ?
              $unsigned(({wire757} ?
                  reg747 : reg739)) : (~&((~^reg755) && $unsigned(reg740)))) ?
          $signed(({wire778[(2'h2):(1'h1)]} < (reg745[(3'h6):(3'h6)] ?
              {reg812,
                  reg695} : ((7'h4a) || reg747)))) : reg730[(1'h1):(1'h0)]))
        begin
          reg816 <= (~^$signed(((~&$signed(reg733)) <= reg783)));
          if ((((8'ha0) ?
                  reg748 : ($signed((reg701 << (8'hba))) ?
                      ({(8'haa)} | $signed(reg781)) : {$signed((8'ha9))})) ?
              (~^$unsigned($unsigned((&reg744)))) : $unsigned(($signed(((7'h41) + reg742)) ?
                  ($unsigned((8'ha2)) ?
                      $unsigned(reg792) : wire766[(1'h0):(1'h0)]) : reg781[(3'h5):(1'h0)]))))
            begin
              reg817 <= reg727[(1'h1):(1'h1)];
              reg818 <= (reg795[(2'h3):(1'h1)] ?
                  reg707 : $signed(reg719[(1'h1):(1'h1)]));
              reg819 <= $signed({reg740,
                  (reg791[(5'h15):(5'h15)] ?
                      (reg705[(2'h2):(2'h2)] ^~ (reg779 == reg696)) : ((reg714 <<< wire692) ?
                          $unsigned(reg790) : ((8'hb6) ^~ (8'ha6))))});
              reg820 <= reg748;
            end
          else
            begin
              reg817 <= (^((reg763[(2'h3):(1'h0)] >= $signed((wire768 ?
                  reg729 : reg769))) - $unsigned(wire775[(3'h5):(1'h1)])));
              reg818 <= ((reg763[(1'h1):(1'h0)] ?
                  reg783[(2'h2):(2'h2)] : $signed((7'h43))) + $signed((|$unsigned($signed(reg726)))));
            end
          reg821 <= $unsigned(((((+reg815) ?
                  ((8'ha6) | reg711) : $unsigned(reg734)) ?
              ($unsigned(reg763) ?
                  (~&reg703) : (reg722 ^ reg709)) : $signed(reg790[(2'h3):(2'h3)])) > ((~^(7'h43)) ?
              ((~|reg724) ?
                  (+reg772) : reg746[(1'h1):(1'h1)]) : ((wire759 & reg792) ?
                  reg735 : (+reg739)))));
          if (reg748[(2'h2):(2'h2)])
            begin
              reg822 <= {reg803,
                  ((($signed(wire690) <= $signed((8'ha3))) ?
                          $unsigned((reg705 ^ reg738)) : $signed($signed(reg781))) ?
                      (reg739[(2'h2):(1'h0)] ?
                          reg788 : ($unsigned(reg714) - (~^reg724))) : reg719[(4'hd):(2'h3)])};
              reg823 <= (^~$signed(reg810[(1'h1):(1'h1)]));
            end
          else
            begin
              reg822 <= (~(({(+(8'ha6)), reg715} ?
                  reg743 : ($unsigned(reg697) ?
                      (reg724 < reg803) : {(8'hbe),
                          wire757})) < (~|((wire759 ^~ reg800) && (wire759 ?
                  reg803 : reg792)))));
              reg823 <= $signed(($signed($signed((wire765 ? reg704 : reg788))) ?
                  (wire767 ?
                      $unsigned(reg747[(2'h2):(1'h0)]) : $unsigned((reg818 ?
                          reg738 : reg703))) : (8'ha1)));
            end
          if ($unsigned($signed($signed(((reg754 ?
              wire761 : reg707) | (!reg724))))))
            begin
              reg824 <= (|(8'hb3));
              reg825 <= $unsigned(reg722[(1'h1):(1'h1)]);
            end
          else
            begin
              reg824 <= $signed(reg780);
              reg825 <= (^~($signed(reg721) ?
                  $signed({$signed(reg771),
                      reg783}) : ($signed(((8'h9c) & reg697)) ?
                      reg751 : (^$unsigned(wire766)))));
              reg826 <= (^~$signed($unsigned({$unsigned(reg813), reg716})));
              reg827 <= $unsigned((&$signed(wire760[(3'h6):(2'h3)])));
              reg828 <= $unsigned(wire759);
            end
        end
      else
        begin
          if ($unsigned({reg718}))
            begin
              reg816 <= (reg755[(3'h5):(3'h4)] ?
                  ($unsigned((reg827[(1'h0):(1'h0)] > {reg720, reg698})) ?
                      ((8'ha2) <= reg763[(2'h2):(2'h2)]) : {(reg741 ?
                              (reg809 >>> reg722) : {reg707}),
                          reg722}) : ($signed(wire765[(4'hc):(4'h8)]) > (($signed(reg805) ?
                      (reg703 - (8'hb2)) : reg751) != reg722[(5'h10):(4'hc)])));
              reg817 <= reg702;
              reg818 <= reg794[(5'h1a):(3'h4)];
            end
          else
            begin
              reg816 <= $unsigned(((reg795[(2'h2):(1'h1)] <= (reg727[(4'h8):(2'h3)] ?
                      $unsigned((8'hb7)) : $signed((8'haf)))) ?
                  reg753 : (({reg803} ?
                          (^wire774) : (reg718 ? reg789 : reg735)) ?
                      reg801[(1'h0):(1'h0)] : $unsigned((8'ha0)))));
              reg817 <= (~$signed(wire778));
              reg818 <= reg784[(3'h7):(2'h3)];
              reg819 <= {$signed(wire776[(2'h3):(2'h2)])};
              reg820 <= (+reg801[(3'h4):(2'h2)]);
              reg821 <= (!$signed($unsigned($signed((&wire777)))));
            end
        end
    end
  assign wire829 = (~$signed(reg824));
  assign wire830 = ((~^$unsigned(reg786[(1'h0):(1'h0)])) + (($unsigned((~|reg710)) ~^ (^(reg763 ?
                       reg712 : reg813))) > $unsigned({$unsigned(reg713)})));
  assign wire831 = (-reg716);
  assign wire832 = $signed(reg817);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module474
#(parameter param633 = (8'h9f))
(y, clk, wire478, wire477, wire476, wire475);
  output wire [(32'h89b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire478;
  input wire [(5'h10):(1'h0)] wire477;
  input wire signed [(5'h10):(1'h0)] wire476;
  input wire signed [(4'hc):(1'h0)] wire475;
  wire signed [(5'h18):(1'h0)] wire632;
  wire [(5'h13):(1'h0)] wire631;
  wire signed [(4'ha):(1'h0)] wire630;
  wire signed [(4'hb):(1'h0)] wire629;
  wire [(4'h9):(1'h0)] wire628;
  wire [(5'h18):(1'h0)] wire627;
  wire [(5'h11):(1'h0)] wire565;
  wire [(2'h2):(1'h0)] wire564;
  wire signed [(5'h11):(1'h0)] wire518;
  wire [(5'h10):(1'h0)] wire494;
  wire signed [(5'h16):(1'h0)] wire493;
  wire signed [(4'hf):(1'h0)] wire492;
  wire signed [(4'hc):(1'h0)] wire491;
  wire [(5'h12):(1'h0)] wire490;
  wire [(5'h15):(1'h0)] wire489;
  wire signed [(4'ha):(1'h0)] wire488;
  wire signed [(4'ha):(1'h0)] wire487;
  wire [(4'ha):(1'h0)] wire486;
  wire [(5'h16):(1'h0)] wire485;
  wire signed [(5'h1a):(1'h0)] wire484;
  wire signed [(3'h5):(1'h0)] wire483;
  wire [(4'hc):(1'h0)] wire482;
  wire [(4'hd):(1'h0)] wire481;
  wire [(5'h12):(1'h0)] wire480;
  wire signed [(4'ha):(1'h0)] wire479;
  reg [(3'h6):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg624 = (1'h0);
  reg [(3'h6):(1'h0)] reg623 = (1'h0);
  reg [(4'he):(1'h0)] reg622 = (1'h0);
  reg [(5'h13):(1'h0)] reg621 = (1'h0);
  reg [(4'hb):(1'h0)] reg620 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg619 = (1'h0);
  reg [(2'h3):(1'h0)] reg618 = (1'h0);
  reg [(3'h7):(1'h0)] reg617 = (1'h0);
  reg [(5'h19):(1'h0)] reg616 = (1'h0);
  reg [(4'h9):(1'h0)] reg615 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg613 = (1'h0);
  reg [(4'hc):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg611 = (1'h0);
  reg [(5'h1a):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg608 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg607 = (1'h0);
  reg [(4'he):(1'h0)] reg606 = (1'h0);
  reg [(5'h16):(1'h0)] reg605 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg604 = (1'h0);
  reg [(4'ha):(1'h0)] reg603 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg601 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg600 = (1'h0);
  reg [(3'h6):(1'h0)] reg599 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg598 = (1'h0);
  reg [(5'h11):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg595 = (1'h0);
  reg [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(3'h4):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg592 = (1'h0);
  reg [(4'h9):(1'h0)] reg591 = (1'h0);
  reg [(3'h7):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg588 = (1'h0);
  reg signed [(4'he):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg585 = (1'h0);
  reg [(4'hc):(1'h0)] reg584 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg582 = (1'h0);
  reg [(5'h1a):(1'h0)] reg581 = (1'h0);
  reg [(4'h9):(1'h0)] reg580 = (1'h0);
  reg [(5'h10):(1'h0)] reg579 = (1'h0);
  reg [(3'h4):(1'h0)] reg578 = (1'h0);
  reg [(5'h12):(1'h0)] reg577 = (1'h0);
  reg [(5'h18):(1'h0)] reg576 = (1'h0);
  reg [(4'he):(1'h0)] reg575 = (1'h0);
  reg [(5'h13):(1'h0)] reg574 = (1'h0);
  reg [(4'h9):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg571 = (1'h0);
  reg [(3'h7):(1'h0)] reg570 = (1'h0);
  reg [(5'h19):(1'h0)] reg569 = (1'h0);
  reg [(5'h12):(1'h0)] reg568 = (1'h0);
  reg [(5'h1a):(1'h0)] reg567 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg566 = (1'h0);
  reg [(2'h2):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg562 = (1'h0);
  reg [(3'h5):(1'h0)] reg561 = (1'h0);
  reg [(2'h2):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg558 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg557 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg556 = (1'h0);
  reg [(5'h19):(1'h0)] reg555 = (1'h0);
  reg [(4'he):(1'h0)] reg554 = (1'h0);
  reg [(3'h7):(1'h0)] reg553 = (1'h0);
  reg [(3'h7):(1'h0)] reg552 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg549 = (1'h0);
  reg [(4'h8):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg546 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg545 = (1'h0);
  reg [(3'h7):(1'h0)] reg544 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg542 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg541 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg540 = (1'h0);
  reg [(5'h13):(1'h0)] reg539 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg537 = (1'h0);
  reg [(4'ha):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg535 = (1'h0);
  reg [(4'h8):(1'h0)] reg534 = (1'h0);
  reg [(2'h2):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg529 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg528 = (1'h0);
  reg [(5'h1a):(1'h0)] reg527 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg526 = (1'h0);
  reg [(3'h6):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg523 = (1'h0);
  reg [(4'ha):(1'h0)] reg522 = (1'h0);
  reg [(4'hb):(1'h0)] reg521 = (1'h0);
  reg [(3'h7):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg519 = (1'h0);
  reg [(5'h17):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg516 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg515 = (1'h0);
  reg [(5'h1a):(1'h0)] reg514 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg513 = (1'h0);
  reg [(5'h11):(1'h0)] reg512 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg509 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg508 = (1'h0);
  reg [(5'h11):(1'h0)] reg507 = (1'h0);
  reg [(5'h11):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg505 = (1'h0);
  reg [(3'h6):(1'h0)] reg504 = (1'h0);
  reg [(4'ha):(1'h0)] reg503 = (1'h0);
  reg [(3'h5):(1'h0)] reg502 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg500 = (1'h0);
  reg [(5'h18):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg498 = (1'h0);
  reg [(5'h14):(1'h0)] reg497 = (1'h0);
  reg [(5'h14):(1'h0)] reg496 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg495 = (1'h0);
  assign y = {wire632,
                 wire631,
                 wire630,
                 wire629,
                 wire628,
                 wire627,
                 wire565,
                 wire564,
                 wire518,
                 wire494,
                 wire493,
                 wire492,
                 wire491,
                 wire490,
                 wire489,
                 wire488,
                 wire487,
                 wire486,
                 wire485,
                 wire484,
                 wire483,
                 wire482,
                 wire481,
                 wire480,
                 wire479,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 (1'h0)};
  assign wire479 = {($unsigned(($signed(wire477) - {wire475})) ?
                           ((wire475 ?
                                   (wire476 > wire478) : (wire478 ?
                                       wire475 : wire477)) ?
                               wire478[(5'h18):(4'hf)] : wire476[(4'hc):(2'h3)]) : wire476[(1'h1):(1'h1)])};
  assign wire480 = wire479;
  assign wire481 = ((($unsigned(((8'hbb) < wire478)) ?
                           (&((8'hb5) ?
                               (8'hb5) : wire478)) : $unsigned({wire475,
                               wire475})) > wire478[(5'h16):(3'h4)]) ?
                       (($signed($unsigned(wire475)) ?
                           wire480 : (wire478[(4'hf):(3'h6)] > wire478)) || $signed($signed((^wire480)))) : wire478[(3'h5):(3'h5)]);
  assign wire482 = (!(($unsigned((8'hb5)) ?
                           (~wire476[(5'h10):(4'hb)]) : ($unsigned((7'h47)) || wire477[(4'ha):(3'h5)])) ?
                       {$signed($signed(wire481)),
                           $unsigned(wire481[(1'h1):(1'h1)])} : wire480));
  assign wire483 = {$unsigned({(^(wire478 ? wire478 : wire480)),
                           $signed($signed(wire476))})};
  assign wire484 = $unsigned(wire475);
  assign wire485 = wire475;
  assign wire486 = wire475;
  assign wire487 = wire486;
  assign wire488 = (wire478[(5'h13):(5'h13)] ?
                       (8'hb6) : wire476[(4'hc):(4'h8)]);
  assign wire489 = (|((wire484[(4'h8):(3'h7)] ?
                           ($signed(wire477) < (&wire483)) : {(wire487 ^~ wire478),
                               $signed(wire481)}) ?
                       wire475[(4'hc):(3'h7)] : (!((wire483 ?
                           wire482 : wire484) - wire485))));
  assign wire490 = $unsigned({{wire477[(3'h4):(1'h0)],
                           (wire485[(5'h15):(5'h12)] ?
                               wire483[(1'h0):(1'h0)] : (wire486 & wire483))}});
  assign wire491 = $signed((^wire479[(4'h8):(3'h4)]));
  assign wire492 = wire489;
  assign wire493 = $unsigned($signed(wire485[(4'h8):(3'h7)]));
  assign wire494 = ($signed((!((wire476 > wire492) + (wire487 ?
                           wire481 : wire486)))) ?
                       (($unsigned($unsigned(wire489)) ?
                           wire483 : $signed(wire480[(5'h12):(4'hd)])) << (8'hba)) : (8'hbc));
  always
    @(posedge clk) begin
      if (wire485[(4'he):(4'h9)])
        begin
          reg495 <= wire488[(2'h2):(2'h2)];
        end
      else
        begin
          reg495 <= $unsigned($signed(wire493));
          if ((~^((~^$signed((~wire490))) >= wire491)))
            begin
              reg496 <= $unsigned($unsigned(wire483[(3'h5):(1'h0)]));
              reg497 <= (7'h4e);
              reg498 <= wire490;
              reg499 <= $unsigned((8'ha9));
              reg500 <= reg496[(4'hb):(3'h4)];
            end
          else
            begin
              reg496 <= ($signed(((~^$unsigned(wire480)) ^ wire482)) ?
                  $unsigned($signed({{wire477,
                          wire480}})) : (({$unsigned(wire477)} ~^ ((wire490 && wire477) ?
                      (8'hbc) : $unsigned(wire485))) < wire476[(1'h1):(1'h0)]));
            end
        end
      if (((8'hac) == $signed(((^~$signed((7'h49))) ?
          ((~&reg497) || $unsigned(wire481)) : $signed($unsigned(reg495))))))
        begin
          if (wire487[(4'h8):(2'h2)])
            begin
              reg501 <= (reg500 | (($unsigned($signed((8'ha4))) << $unsigned($unsigned((7'h4e)))) ?
                  (8'ha8) : $signed($signed(wire478[(4'hc):(2'h2)]))));
              reg502 <= (+{$signed($unsigned($unsigned(wire479))),
                  $signed((-(wire494 ? (8'h9e) : (7'h45))))});
            end
          else
            begin
              reg501 <= $signed(wire483);
              reg502 <= (((((-wire483) ?
                  (wire479 >> wire481) : $unsigned(reg499)) == $unsigned(((8'ha6) ~^ reg498))) <<< (^(&wire489))) & $unsigned((((reg497 >= wire481) <= (wire478 ?
                  wire477 : reg500)) ^~ wire492[(3'h6):(2'h3)])));
              reg503 <= (^~$signed((wire487 < {$signed(wire493),
                  $signed(wire491)})));
            end
          reg504 <= $unsigned({(wire493 ?
                  $signed((reg499 ? reg500 : wire489)) : $unsigned(wire480)),
              {$unsigned((wire487 <= reg503)), wire492[(4'h8):(4'h8)]}});
          if ({reg496,
              ((!(&wire488[(3'h6):(1'h0)])) ?
                  (+(8'hbb)) : (reg504 ?
                      $unsigned({reg497, reg500}) : {wire483}))})
            begin
              reg505 <= $signed(reg500);
              reg506 <= $signed((7'h43));
              reg507 <= wire484;
              reg508 <= {(($unsigned((~reg495)) ?
                      wire494 : (-reg496)) <= $signed((~(reg504 ^ wire493)))),
                  $unsigned((((wire484 < wire484) - $signed(reg499)) ?
                      wire483 : (~&$unsigned((8'hbf)))))};
            end
          else
            begin
              reg505 <= $signed($unsigned(((^(wire486 & (8'h9e))) >= ($unsigned(wire493) | $unsigned(wire477)))));
              reg506 <= $signed((wire492[(4'hd):(2'h3)] ~^ reg499[(4'hc):(3'h6)]));
              reg507 <= $signed($unsigned($unsigned(((^~reg495) ?
                  $signed(wire484) : (~^wire485)))));
              reg508 <= wire483[(1'h1):(1'h1)];
              reg509 <= wire477[(4'h8):(4'h8)];
              reg510 <= (~|$signed(wire490));
            end
          if ($unsigned((8'hb6)))
            begin
              reg511 <= (|$signed((-(reg504 <= $unsigned(reg509)))));
              reg512 <= {({$signed((wire485 ? (8'hb5) : wire476))} ?
                      $signed(reg506[(4'he):(4'hb)]) : $signed(((reg511 ^~ wire477) ?
                          ((8'hb7) ? reg505 : reg499) : (wire482 == wire485)))),
                  {reg497}};
              reg513 <= (((~|wire489[(5'h14):(5'h13)]) ?
                      wire484[(4'h9):(3'h6)] : {reg500[(4'hd):(1'h0)],
                          (reg502 ~^ (~&reg503))}) ?
                  wire494[(4'h8):(1'h0)] : wire488[(3'h4):(2'h2)]);
              reg514 <= (&$signed(wire482));
              reg515 <= $signed((((~&$signed(wire488)) ~^ $unsigned(wire483)) ?
                  (reg498 ?
                      wire481[(4'ha):(1'h0)] : $unsigned((wire484 ?
                          wire483 : (8'hb1)))) : $unsigned(($unsigned((8'hb3)) ?
                      $signed(wire493) : (7'h4b)))));
              reg516 <= $unsigned({(8'ha1),
                  {{(reg499 ? reg496 : wire479), $signed(wire493)},
                      $signed($unsigned(reg513))}});
            end
          else
            begin
              reg511 <= $unsigned($signed(wire490));
              reg512 <= ((($signed($unsigned(reg501)) ?
                      (reg495 & $unsigned(reg510)) : reg511) ?
                  $unsigned($signed($signed(wire494))) : (($signed((8'haa)) ~^ wire483[(2'h2):(1'h1)]) + wire494[(4'ha):(1'h1)])) << wire477[(3'h5):(3'h4)]);
              reg513 <= reg499;
              reg514 <= (|$signed($unsigned(wire481)));
            end
          reg517 <= $unsigned((wire479[(4'h9):(3'h6)] ?
              $unsigned(reg498[(1'h1):(1'h1)]) : $unsigned((7'h4e))));
        end
      else
        begin
          if (wire492[(2'h3):(2'h2)])
            begin
              reg501 <= $signed(reg498[(3'h5):(1'h1)]);
              reg502 <= wire480[(4'hf):(3'h4)];
            end
          else
            begin
              reg501 <= $signed((&$unsigned((~&(reg507 <= (8'hac))))));
              reg502 <= {((~&wire482) ?
                      {({(7'h45), reg499} ?
                              wire494 : $signed(reg510))} : (8'hb0)),
                  wire490[(3'h5):(2'h3)]};
              reg503 <= $signed($signed($signed($unsigned((reg513 >>> reg513)))));
            end
          if (wire480)
            begin
              reg504 <= {{{(~|wire487[(2'h2):(1'h0)]), (~$signed(reg498))}},
                  ((|(((7'h4d) ? wire488 : reg503) && (reg501 ?
                      reg497 : reg515))) <= ($signed(reg497[(4'h9):(3'h6)]) << ($signed((8'hb0)) - ((8'had) ?
                      reg505 : wire480))))};
              reg505 <= $unsigned($signed({wire481}));
              reg506 <= (^~(7'h44));
              reg507 <= (|($unsigned($unsigned(reg499[(5'h11):(2'h3)])) ^ $signed((wire491[(3'h4):(2'h3)] ?
                  $unsigned(wire480) : (wire476 != reg511)))));
              reg508 <= reg506[(3'h6):(3'h5)];
            end
          else
            begin
              reg504 <= $unsigned({(+((reg517 ? wire477 : reg501) ^ {wire493})),
                  (reg512 ? reg495 : wire480[(4'he):(3'h6)])});
              reg505 <= $unsigned(((reg499[(3'h5):(3'h4)] < ((reg511 ?
                      wire487 : (7'h4b)) ?
                  wire483[(1'h1):(1'h0)] : wire488[(4'h8):(3'h7)])) ^~ $unsigned((wire479 - $signed(wire475)))));
              reg506 <= $signed(((|wire482) ?
                  $signed({(reg497 ? (8'hab) : (8'hb7)),
                      (|wire476)}) : $signed($unsigned((~&(8'hb6))))));
              reg507 <= ($unsigned(wire494) ? (~wire488) : wire480);
              reg508 <= (!{reg503, $unsigned(reg497)});
            end
          reg509 <= {$unsigned({reg506, (wire487 & wire492[(3'h6):(3'h4)])}),
              ($signed((reg514[(5'h16):(4'ha)] ^ (wire479 ?
                  reg514 : reg497))) + ($signed({reg504}) + ((&wire493) <= reg507)))};
        end
    end
  assign wire518 = ($unsigned($signed((7'h46))) ?
                       ((~&$unsigned($signed(reg510))) ?
                           {$unsigned((+reg503))} : (($signed(reg515) > $unsigned((7'h40))) << $unsigned({reg514}))) : (($unsigned((wire492 ?
                                   wire478 : wire493)) ?
                               $signed(reg502[(2'h3):(2'h2)]) : (~|{reg506,
                                   wire492})) ?
                           (&(&wire477)) : $signed((8'ha2))));
  always
    @(posedge clk) begin
      if ((($signed(wire481) ?
              wire479 : (reg502 >= $signed($unsigned(wire491)))) ?
          (((~&wire488) ~^ wire483) ^~ $unsigned((&$signed(reg511)))) : wire479[(3'h6):(3'h6)]))
        begin
          reg519 <= (^reg516);
          reg520 <= $unsigned(($signed($unsigned(wire493[(4'ha):(3'h7)])) ?
              $unsigned({{wire475},
                  $unsigned(reg516)}) : (reg509[(3'h6):(3'h4)] ?
                  (reg502[(3'h4):(2'h2)] ?
                      (reg515 ?
                          reg499 : reg502) : (reg510 > reg501)) : reg515)));
        end
      else
        begin
          reg519 <= $unsigned((wire479 ?
              (($unsigned(reg512) ? reg515 : (reg497 ? reg501 : wire475)) ?
                  ($signed(reg509) ?
                      wire493 : wire488) : (~|wire486)) : (~&$signed((wire491 ?
                  reg514 : (8'ha9))))));
        end
      reg521 <= $signed((^~(!($signed(wire488) + (wire491 ?
          wire490 : wire489)))));
      reg522 <= ({wire479[(4'ha):(2'h2)], $unsigned(reg509)} ?
          reg507 : $signed((+(^~wire481[(3'h4):(3'h4)]))));
      if (wire489)
        begin
          if (wire485)
            begin
              reg523 <= $unsigned((&((!(wire485 == reg510)) ?
                  {(wire482 > reg521)} : ($unsigned((8'h9f)) ?
                      wire486 : reg504[(3'h6):(1'h1)]))));
              reg524 <= {(wire493[(5'h12):(4'h9)] <= (((~|wire482) - reg502[(3'h4):(1'h1)]) ^ {(wire483 < reg509),
                      wire482[(4'hc):(3'h5)]}))};
              reg525 <= ($signed((&reg516)) ?
                  reg506 : $unsigned({(reg511 | (^~wire489)),
                      (~^{reg521, wire476})}));
              reg526 <= reg515;
              reg527 <= wire486;
            end
          else
            begin
              reg523 <= reg516[(4'ha):(3'h6)];
              reg524 <= wire489[(4'ha):(1'h0)];
              reg525 <= reg508;
              reg526 <= $signed($signed(($unsigned((^~(7'h43))) ?
                  ({wire480, wire494} ?
                      reg513[(2'h2):(1'h1)] : {reg519}) : ((~^(8'h9f)) <<< reg512[(4'he):(4'he)]))));
              reg527 <= $unsigned($signed($signed(reg517)));
              reg528 <= ((reg519[(3'h5):(3'h5)] | (-(!(wire475 && wire493)))) ?
                  (^~reg525) : {$signed($signed($signed(reg495)))});
            end
          if ((~|(((wire493 ? $signed((8'hbb)) : (reg506 ^ reg528)) ?
              $unsigned((reg499 ?
                  reg520 : reg508)) : $unsigned((^(8'hb5)))) ~^ wire486[(3'h4):(2'h2)])))
            begin
              reg529 <= ((!(((reg528 - reg497) ?
                  (8'hab) : $signed(reg510)) << $unsigned($signed(wire486)))) < $signed(($unsigned((wire488 ?
                      wire484 : reg514)) ?
                  ($signed(reg500) * (reg510 ? reg495 : reg502)) : ((wire518 ?
                          wire518 : (8'h9f)) ?
                      $unsigned(wire490) : (wire518 ^~ (8'hb2))))));
              reg530 <= {(({(wire478 ? reg514 : (8'haa)), $unsigned(reg505)} ?
                          reg510 : reg510) ?
                      wire492[(3'h7):(2'h2)] : (wire477[(2'h2):(2'h2)] ?
                          $unsigned((wire491 ?
                              (7'h45) : reg513)) : ((wire491 ^~ reg502) << (reg496 < reg506)))),
                  (~|(reg521[(4'hb):(3'h7)] >= (wire492 > reg496[(3'h6):(1'h0)])))};
              reg531 <= wire487;
              reg532 <= {$unsigned({reg511[(3'h6):(2'h2)]}),
                  reg508[(3'h7):(3'h7)]};
              reg533 <= $unsigned({reg514, $signed((^(wire486 != wire488)))});
            end
          else
            begin
              reg529 <= reg495[(2'h3):(1'h0)];
              reg530 <= $signed($signed((~^$signed(reg520))));
              reg531 <= reg530;
            end
          reg534 <= (wire485[(4'h9):(3'h6)] ^ (!wire518[(3'h6):(3'h5)]));
          reg535 <= wire490;
          if ((-(~|({reg515[(2'h2):(1'h1)]} | (wire480 ?
              $signed((7'h4b)) : $signed(reg525))))))
            begin
              reg536 <= reg517[(5'h15):(3'h7)];
              reg537 <= (8'hba);
              reg538 <= $unsigned((~^wire476[(4'hf):(1'h0)]));
              reg539 <= $signed(reg507);
              reg540 <= (!$unsigned(($signed((-wire477)) <<< (!$unsigned((8'hb7))))));
              reg541 <= $unsigned(reg536);
            end
          else
            begin
              reg536 <= wire478[(3'h7):(3'h6)];
              reg537 <= $unsigned(((reg514[(5'h15):(4'hb)] ?
                  reg506[(3'h7):(3'h5)] : ($signed(wire493) ?
                      reg515[(2'h3):(2'h2)] : $signed(reg506))) && (((8'hbb) ?
                      (wire481 ? wire475 : (8'hb5)) : reg538[(4'h9):(1'h1)]) ?
                  $unsigned(reg541[(4'hb):(1'h0)]) : (~$unsigned(reg505)))));
              reg538 <= (wire491 ?
                  $unsigned(((wire479[(3'h7):(3'h4)] ?
                          (~|reg505) : reg510[(5'h10):(4'hb)]) ?
                      wire492 : (^(wire483 ?
                          wire489 : reg507)))) : $signed($signed($unsigned($signed(wire481)))));
              reg539 <= (^$signed(wire484));
            end
          if ($unsigned(wire482[(2'h2):(2'h2)]))
            begin
              reg542 <= $signed($unsigned(((8'hb2) ?
                  ($signed(wire479) ?
                      (reg507 ?
                          reg510 : reg529) : reg519[(4'h9):(3'h5)]) : $signed((+reg503)))));
              reg543 <= (wire488[(2'h3):(1'h0)] ?
                  $unsigned(reg511[(4'h9):(3'h5)]) : $unsigned($unsigned(wire481[(2'h3):(1'h1)])));
              reg544 <= (+reg502);
              reg545 <= ($signed(reg530[(5'h14):(1'h0)]) ?
                  ((|(&reg511)) ?
                      wire492 : $unsigned(reg500[(4'ha):(3'h4)])) : $unsigned((&$signed($signed(reg506)))));
              reg546 <= {{$signed((8'h9d))},
                  $unsigned($signed($signed(reg526[(1'h1):(1'h1)])))};
            end
          else
            begin
              reg542 <= (8'hb2);
              reg543 <= reg495;
              reg544 <= (reg542[(5'h12):(5'h10)] >= $signed((((-reg524) <= {(8'h9c),
                  reg541}) != wire488)));
              reg545 <= reg546;
              reg546 <= reg522;
            end
        end
      else
        begin
          reg523 <= (|wire488);
          reg524 <= {$unsigned((({reg524} ?
                      (wire476 ? (8'hb6) : (8'hab)) : (wire493 ~^ reg521)) ?
                  $signed(reg505) : $signed(reg525))),
              {reg542[(3'h4):(3'h4)],
                  (-((^(8'hba)) ~^ reg508[(3'h6):(3'h5)]))}};
        end
      if (($signed(reg528) >= reg526))
        begin
          if (($signed((($signed(reg497) <<< (wire490 ? reg529 : reg511)) ?
              $unsigned(reg509[(4'hf):(3'h7)]) : $unsigned($signed(reg514)))) < (~^(^~(|$unsigned(wire480))))))
            begin
              reg547 <= ($unsigned((((wire481 ? reg516 : reg505) ?
                          reg506[(3'h6):(1'h0)] : $unsigned((8'ha5))) ?
                      ({wire518, reg498} ?
                          (!wire484) : $unsigned((8'hb0))) : reg519[(4'hd):(4'h8)])) ?
                  ($signed(reg509) + reg500) : (~^reg525));
            end
          else
            begin
              reg547 <= $signed($unsigned((((reg507 ?
                      reg533 : wire475) ^ (reg535 + reg533)) ?
                  reg541[(3'h4):(1'h1)] : ($signed(reg545) ?
                      (reg513 ? wire487 : reg505) : reg514))));
            end
          reg548 <= $unsigned(reg540[(1'h1):(1'h0)]);
        end
      else
        begin
          reg547 <= (((~^{$unsigned(reg527),
              (reg509 ? wire487 : reg511)}) + (reg525 ?
              $signed($unsigned(reg521)) : (~&(!(7'h40))))) <= reg498);
          reg548 <= (!(reg496 && $unsigned($unsigned({reg510}))));
          reg549 <= wire489[(1'h0):(1'h0)];
          reg550 <= (reg544 >> $signed(reg506[(2'h2):(2'h2)]));
          if ($signed(((^(reg499 >> $unsigned(reg550))) ?
              $signed(((wire487 >= reg523) ?
                  (reg538 ?
                      wire489 : (8'hb8)) : $unsigned(reg524))) : $signed((~&(reg524 ?
                  reg549 : reg550))))))
            begin
              reg551 <= $signed((~{($signed(reg514) ?
                      {wire490, (8'ha7)} : $unsigned(reg539))}));
            end
          else
            begin
              reg551 <= reg502[(2'h3):(2'h2)];
              reg552 <= wire518;
              reg553 <= $signed((^reg506));
              reg554 <= $signed(wire491[(3'h4):(2'h3)]);
              reg555 <= $signed(reg502[(2'h3):(1'h1)]);
              reg556 <= $signed((8'hae));
            end
          if ($unsigned(wire487))
            begin
              reg557 <= $unsigned($unsigned(reg533));
              reg558 <= {reg522, reg555[(1'h0):(1'h0)]};
              reg559 <= reg558[(4'h8):(3'h7)];
              reg560 <= $signed($signed(((8'ha8) ?
                  reg554[(3'h4):(2'h2)] : $unsigned(wire480))));
            end
          else
            begin
              reg557 <= reg560[(1'h1):(1'h1)];
              reg558 <= wire482;
              reg559 <= $unsigned(wire482);
              reg560 <= (^(($unsigned((reg531 || reg512)) - reg526) * (8'h9f)));
              reg561 <= $unsigned(reg501);
              reg562 <= $unsigned(($unsigned(($signed(reg520) >= $signed(reg517))) ?
                  $unsigned({$signed((7'h4a))}) : (reg505 ~^ ((reg549 * reg533) + $unsigned(wire481)))));
            end
        end
      reg563 <= (({$unsigned($signed(reg554))} ?
              (reg557 == reg527) : {(7'h4b), $unsigned((reg552 != reg549))}) ?
          wire481 : reg552[(3'h5):(3'h4)]);
    end
  assign wire564 = $signed(reg540[(2'h3):(2'h2)]);
  assign wire565 = (~reg506);
  always
    @(posedge clk) begin
      if (({(8'hb9)} ?
          ((-(!{reg505})) >> (reg532[(3'h4):(3'h4)] ?
              (~|reg503) : reg514)) : (reg505 ?
              $unsigned($signed((8'ha6))) : (~&((reg527 ? reg554 : (8'hab)) ?
                  reg509[(4'hf):(4'he)] : $signed(reg536))))))
        begin
          if ((^(reg515[(3'h5):(1'h0)] ^ $signed($signed((8'hb6))))))
            begin
              reg566 <= ($unsigned(($signed((^reg521)) >= (~&wire565))) ^ ((($signed(reg542) ^~ $signed((8'h9d))) <<< ($unsigned((8'hb4)) ?
                      (reg524 ? (8'h9c) : wire476) : (reg561 > wire476))) ?
                  {{wire482,
                          reg537}} : $signed($signed(((8'ha7) >= (8'hab))))));
              reg567 <= (^$unsigned($signed((reg539[(3'h6):(1'h1)] ?
                  (reg555 > reg528) : (&reg542)))));
              reg568 <= (^~(|$signed(($unsigned(reg531) ?
                  (~(8'ha2)) : (-reg495)))));
              reg569 <= {$signed(reg495[(1'h1):(1'h0)]),
                  $signed(wire492[(4'he):(3'h5)])};
            end
          else
            begin
              reg566 <= (~|(!$signed(wire493)));
              reg567 <= (($signed($signed(reg510[(4'he):(1'h0)])) ?
                  $unsigned(reg555) : reg521) ^ reg527[(5'h12):(4'h9)]);
            end
          if (reg556[(1'h0):(1'h0)])
            begin
              reg570 <= reg497;
              reg571 <= reg539;
            end
          else
            begin
              reg570 <= $unsigned($signed((!reg496)));
              reg571 <= {($signed({(reg544 ? reg532 : (8'ha8)),
                      reg532[(4'h9):(3'h6)]}) > ((reg529[(4'he):(4'ha)] ?
                      (reg497 < wire480) : reg525[(2'h2):(2'h2)]) <<< ((wire488 ?
                          (8'hb2) : reg562) ?
                      (~|reg529) : {wire491, reg544}))),
                  {(7'h48)}};
              reg572 <= $signed((wire482[(1'h0):(1'h0)] <= reg527));
              reg573 <= (-(^~$signed(wire484[(4'he):(3'h6)])));
              reg574 <= (^~$signed(($signed($unsigned(reg553)) ?
                  $signed($unsigned(wire486)) : $signed($unsigned(wire483)))));
            end
          if (wire494[(4'hf):(4'hb)])
            begin
              reg575 <= reg544;
              reg576 <= $signed(($signed(wire484[(4'hf):(3'h5)]) ?
                  {(reg569[(5'h17):(4'hb)] >= (reg523 || reg509))} : ((reg562[(1'h1):(1'h0)] ?
                      wire490 : {reg536, reg523}) * (+(reg511 ?
                      reg550 : reg540)))));
            end
          else
            begin
              reg575 <= $signed(((reg529[(5'h13):(4'he)] ?
                  {((7'h4b) ?
                          reg504 : reg549)} : (~(!wire565))) | ((~&$signed(reg529)) ?
                  (~|$signed(wire475)) : $unsigned((|reg555)))));
              reg576 <= {(((8'hb2) ?
                          (-(wire564 ? wire479 : wire480)) : ($signed(wire484) ?
                              (~wire565) : $unsigned(reg515))) ?
                      {(reg544[(2'h3):(1'h0)] ?
                              (~reg534) : $unsigned(reg501))} : (8'hb4))};
              reg577 <= reg572;
              reg578 <= (8'ha4);
            end
          if (reg550[(3'h6):(2'h2)])
            begin
              reg579 <= (8'hbb);
              reg580 <= reg503;
              reg581 <= $signed($signed((~|reg501)));
              reg582 <= $signed($signed((~($signed(reg574) <= {(8'ha6),
                  wire477}))));
            end
          else
            begin
              reg579 <= $signed($signed($signed(reg545)));
              reg580 <= (8'hbb);
              reg581 <= reg515[(3'h5):(1'h1)];
              reg582 <= (reg568 == $unsigned($signed({(reg523 ?
                      reg568 : reg562),
                  (reg500 == (8'haa))})));
              reg583 <= $signed(reg561[(2'h2):(1'h1)]);
              reg584 <= ($unsigned(wire490) ^~ reg568);
            end
        end
      else
        begin
          reg566 <= (reg579 ?
              (&(wire489 <= {(reg503 * reg528),
                  (~reg527)})) : wire484[(4'ha):(2'h3)]);
          reg567 <= $signed(reg503[(1'h0):(1'h0)]);
          if ($unsigned(((reg502 - ((wire483 == wire492) ^ (reg542 != reg501))) >>> wire492[(4'hd):(3'h7)])))
            begin
              reg568 <= reg577[(4'hc):(4'h8)];
              reg569 <= $unsigned(reg530[(4'hc):(4'hc)]);
              reg570 <= ($unsigned($unsigned($signed($unsigned((8'had))))) & $signed(((&(reg521 ?
                      reg533 : wire487)) ?
                  (reg577 > (reg550 - reg558)) : (^$signed(reg562)))));
              reg571 <= ($signed((!$signed(reg501[(2'h2):(2'h2)]))) ?
                  (reg571 ?
                      reg520[(3'h6):(1'h0)] : $unsigned(((8'h9e) != (reg526 > (7'h45))))) : {$signed({reg581,
                          reg523})});
            end
          else
            begin
              reg568 <= ((((reg524 ?
                      reg528[(3'h4):(1'h1)] : {reg512}) && reg580) ?
                  $unsigned($signed((reg582 ?
                      wire477 : (8'ha2)))) : (|$unsigned(reg513[(4'hf):(3'h5)]))) >> wire479);
              reg569 <= wire482[(1'h1):(1'h1)];
              reg570 <= {$signed($signed($unsigned((reg501 ?
                      reg524 : reg538)))),
                  (($signed($unsigned(reg501)) * reg508) + (reg562 ?
                      ((reg569 * wire492) ?
                          (reg544 ? reg535 : reg505) : (reg555 ?
                              reg582 : reg584)) : reg566))};
              reg571 <= ($signed(reg511[(4'h8):(1'h1)]) ~^ (^($unsigned({reg568,
                      reg549}) ?
                  (-$signed(reg543)) : $unsigned(reg527[(5'h19):(5'h14)]))));
              reg572 <= ((~|$signed(reg502)) ?
                  ($signed(((~|(7'h42)) ?
                          reg536[(4'ha):(4'h8)] : (reg547 && reg570))) ?
                      $unsigned(reg542) : {(~^(reg498 == (8'ha5)))}) : $unsigned(wire482));
            end
        end
      if (({reg497[(4'h9):(1'h1)]} != (8'h9e)))
        begin
          reg585 <= (+reg551[(3'h5):(1'h1)]);
          reg586 <= reg571[(5'h10):(4'hd)];
          reg587 <= reg558[(4'he):(1'h1)];
        end
      else
        begin
          if ($signed(reg541[(3'h6):(2'h3)]))
            begin
              reg585 <= reg578;
              reg586 <= {$signed($signed($unsigned($signed(reg553))))};
            end
          else
            begin
              reg585 <= $signed((!{$signed($signed(wire491)),
                  {(reg545 ? reg562 : wire486)}}));
              reg586 <= $signed((wire488 <= (((^reg541) ?
                  (reg557 ?
                      wire476 : reg501) : $unsigned(reg567)) * $unsigned(reg580[(3'h5):(1'h0)]))));
              reg587 <= (reg571 > $unsigned($unsigned(reg515)));
              reg588 <= ((~|($unsigned((wire487 ?
                      reg557 : reg566)) > $signed((reg527 ?
                      reg579 : wire482)))) ?
                  reg550[(1'h0):(1'h0)] : {(reg551[(1'h0):(1'h0)] ?
                          ((reg548 > wire485) ?
                              (wire477 ? reg554 : reg571) : (reg551 ?
                                  reg579 : reg500)) : $signed((wire490 ?
                              wire494 : reg581))),
                      $unsigned(($unsigned((8'hb3)) ?
                          $unsigned((8'hb8)) : (reg532 ~^ reg578)))});
              reg589 <= (|((reg504 ?
                      ($unsigned(reg567) ?
                          reg544 : reg566) : reg569[(3'h4):(2'h2)]) ?
                  ($signed((!reg502)) ?
                      (!(reg533 ?
                          wire565 : reg577)) : $unsigned((reg524 | (8'hb4)))) : reg570[(3'h7):(3'h4)]));
              reg590 <= (reg515 << (^~$unsigned((reg502 < reg527[(5'h16):(5'h14)]))));
            end
          reg591 <= reg510;
          reg592 <= $signed($unsigned(reg501[(4'he):(4'h9)]));
          if ((($signed(((reg538 >>> (8'hbe)) || $unsigned(reg504))) <= ($unsigned(reg559) ?
                  reg533 : reg561)) ?
              reg560[(2'h2):(1'h1)] : (~|(((reg505 ?
                  reg590 : reg549) >= ((7'h4b) == (7'h4d))) >= $signed($signed((8'h9c)))))))
            begin
              reg593 <= reg514[(2'h2):(1'h1)];
              reg594 <= (((^~$signed((~&(8'hb4)))) >>> reg498[(3'h6):(3'h5)]) == {(^$unsigned($unsigned(reg515)))});
              reg595 <= {reg517[(2'h3):(2'h3)], (-wire480[(3'h7):(3'h4)])};
              reg596 <= wire489;
              reg597 <= (~&{$signed($signed($signed(reg578)))});
              reg598 <= $signed((wire481 ?
                  (((!(8'ha9)) ? (reg529 >> reg537) : (reg496 + (8'hbb))) ?
                      $signed(reg581[(5'h1a):(4'hf)]) : wire477[(4'he):(3'h5)]) : (~&{(!reg509)})));
            end
          else
            begin
              reg593 <= reg502[(1'h1):(1'h1)];
              reg594 <= $signed(reg548[(4'h8):(2'h2)]);
              reg595 <= (-reg544[(3'h4):(2'h3)]);
              reg596 <= (((+(reg516 ?
                      (-reg589) : $unsigned(reg571))) - wire564) ?
                  ($signed(reg589) ?
                      (+reg563[(1'h1):(1'h0)]) : ($unsigned(((7'h40) ?
                              reg513 : reg586)) ?
                          ({reg516, wire485} ?
                              (reg550 ?
                                  (8'hbf) : wire491) : $signed(reg527)) : $unsigned((reg570 ?
                              reg595 : reg519)))) : $unsigned($unsigned((!((8'hb2) ~^ (8'hba))))));
            end
          if ({(reg554 ? reg535[(2'h2):(1'h1)] : reg505[(1'h1):(1'h1)])})
            begin
              reg599 <= wire486;
              reg600 <= $unsigned((~^({$signed(reg599), (reg525 <= reg590)} ?
                  ($signed(reg498) == (reg553 ?
                      (8'h9e) : reg503)) : reg497[(2'h2):(2'h2)])));
              reg601 <= (reg508[(1'h1):(1'h0)] ?
                  ((|$signed((reg591 >= reg496))) ?
                      {$signed(reg567[(5'h1a):(5'h13)]),
                          wire485} : (8'h9f)) : $signed($signed({(~|reg537),
                      reg526})));
              reg602 <= ($unsigned((~&$unsigned(reg543[(2'h2):(1'h1)]))) ?
                  (($signed({reg522}) ~^ $signed((!reg497))) ^~ ((|(reg498 >= wire493)) ?
                      reg523[(5'h11):(4'hd)] : $unsigned(reg547))) : (((-reg551) ?
                      (^wire564[(1'h1):(1'h0)]) : reg583[(2'h3):(2'h3)]) > reg537[(5'h14):(2'h3)]));
            end
          else
            begin
              reg599 <= (wire483 || reg537);
              reg600 <= {(reg503 ?
                      reg600[(2'h2):(1'h0)] : reg581[(1'h1):(1'h1)]),
                  (reg559[(2'h2):(1'h1)] != reg586)};
              reg601 <= (reg590[(2'h2):(1'h1)] ?
                  ($signed((8'hab)) * $unsigned(($signed((8'h9d)) < ((8'hb0) ?
                      reg602 : reg566)))) : ($unsigned({reg566,
                      $unsigned(wire480)}) ^ $signed(((reg573 * reg527) ^~ ((8'hae) >> reg538)))));
              reg602 <= {(($unsigned((reg568 ? wire491 : (8'h9d))) ?
                      ((+reg595) ?
                          reg543[(3'h5):(2'h3)] : reg531[(5'h16):(4'hd)]) : $unsigned((reg522 < reg531))) == reg549),
                  (&($unsigned({reg553, (8'hab)}) ?
                      (((7'h4e) ? (8'hbc) : reg495) ?
                          (|reg510) : (|reg506)) : $unsigned((|reg554))))};
            end
        end
      reg603 <= (-$signed($unsigned(reg522[(3'h6):(1'h1)])));
      if ((wire482 ?
          {(((reg566 ? (8'hbe) : reg577) ^~ $unsigned((8'hb2))) ?
                  {(reg572 ? reg597 : reg501)} : {(wire482 ?
                          (7'h47) : wire483)}),
              (reg556 - reg522[(3'h6):(2'h2)])} : (({reg592} ?
                  $signed($unsigned(reg527)) : reg528) ?
              (($unsigned(reg519) >>> (wire476 ? reg547 : reg585)) ?
                  ((reg535 * reg603) ?
                      (reg529 ? reg525 : reg498) : (reg502 ?
                          reg584 : (8'had))) : (!(reg566 ?
                      wire482 : reg560))) : (((reg545 ~^ reg584) < (7'h4c)) << $unsigned((-(8'hb3)))))))
        begin
          reg604 <= (&wire486);
          if ((~^$unsigned(($unsigned($unsigned((7'h46))) ?
              (7'h4e) : $unsigned($unsigned(wire564))))))
            begin
              reg605 <= (~reg571);
              reg606 <= (reg569 ? reg506 : $unsigned(reg580));
              reg607 <= (wire478[(4'h8):(1'h1)] ?
                  $unsigned((wire480 ?
                      reg585[(3'h7):(3'h7)] : ($signed((8'hb8)) < reg586[(4'hd):(3'h4)]))) : reg536[(3'h6):(3'h5)]);
            end
          else
            begin
              reg605 <= reg551[(3'h5):(2'h3)];
              reg606 <= reg605[(5'h10):(4'he)];
              reg607 <= (8'haf);
              reg608 <= (reg571[(5'h12):(5'h11)] & ($unsigned(reg566) && ((|{wire478}) * reg510)));
              reg609 <= $signed($signed((($unsigned(reg563) ?
                      $unsigned(reg533) : {reg591}) ?
                  $signed((reg532 ? wire564 : reg540)) : {(reg606 < reg511)})));
            end
          if ($signed(((((reg507 ? reg602 : wire489) | (wire492 ?
                  reg596 : reg526)) != reg495) ?
              $unsigned(($unsigned(wire491) ?
                  (reg499 < reg514) : reg558[(3'h5):(1'h0)])) : (7'h42))))
            begin
              reg610 <= $unsigned(((($signed(reg503) > (reg527 ?
                  reg598 : reg591)) >= wire494[(4'hb):(4'h8)]) != (+$unsigned($unsigned(reg519)))));
              reg611 <= (({reg576[(3'h6):(2'h2)],
                          $unsigned($unsigned(reg581))} ?
                      ({(reg603 | reg509)} ?
                          ((^reg499) ?
                              $signed(reg534) : wire493[(4'hf):(3'h6)]) : $signed((!reg504))) : reg588) ?
                  ({((^reg559) ~^ (reg547 ? reg538 : reg496)),
                          ($unsigned(reg526) ~^ (|(8'hbb)))} ?
                      (((reg549 & reg568) ? $signed((8'ha5)) : (|(7'h43))) ?
                          (~((8'ha0) ? wire475 : (8'ha6))) : ((reg523 ?
                              reg549 : reg548) <= wire564)) : reg598) : (($signed({reg562}) ?
                      reg576[(2'h3):(2'h2)] : (-wire492)) > reg552));
              reg612 <= $signed(((+($signed((8'hb3)) ?
                  $unsigned(reg535) : (reg501 > reg601))) > {(|wire487[(4'h9):(4'h8)])}));
              reg613 <= (8'ha1);
              reg614 <= reg588;
            end
          else
            begin
              reg610 <= $signed(reg536);
              reg611 <= $signed($unsigned(wire481[(4'hd):(4'ha)]));
              reg612 <= $unsigned(wire493);
              reg613 <= $signed(((reg517 != reg498) ?
                  wire476 : reg534[(4'h8):(3'h7)]));
              reg614 <= $signed($signed($signed(reg596[(4'h8):(3'h6)])));
            end
        end
      else
        begin
          if (({$unsigned($signed(wire484)),
              $signed(reg577)} > (reg531 & $unsigned(reg611[(5'h10):(1'h0)]))))
            begin
              reg604 <= (({$signed(reg495), $signed($unsigned((8'h9e)))} ?
                  $signed(($signed(reg537) ^ ((8'ha9) != reg580))) : $signed((~|$unsigned(reg512)))) >= (~&$signed($signed($signed(wire478)))));
              reg605 <= ($signed(wire483[(2'h3):(1'h1)]) <<< $unsigned(reg604[(2'h3):(1'h1)]));
              reg606 <= $signed((reg510 <<< ($signed((^~reg595)) ?
                  $signed({reg507}) : (reg573[(3'h4):(3'h4)] ?
                      (&reg530) : wire494))));
              reg607 <= reg548[(2'h3):(1'h0)];
            end
          else
            begin
              reg604 <= $signed($signed($signed($unsigned($unsigned(reg607)))));
              reg605 <= reg607[(2'h2):(1'h1)];
            end
          reg608 <= $signed(reg527[(5'h15):(4'h9)]);
        end
      if ((($unsigned(reg499) <= $unsigned((&(^reg553)))) == $unsigned(reg553[(1'h0):(1'h0)])))
        begin
          reg615 <= reg605[(3'h5):(1'h0)];
        end
      else
        begin
          if ((reg536 ?
              $unsigned((reg519[(2'h2):(1'h0)] ?
                  {(|(8'haf)),
                      $signed(reg572)} : {reg552[(1'h0):(1'h0)]})) : (~|$signed(reg590[(3'h5):(1'h1)]))))
            begin
              reg615 <= $unsigned($signed($unsigned((^~reg589))));
              reg616 <= ($signed($signed((reg511 & ((8'hae) ^ reg549)))) || (7'h49));
              reg617 <= $signed($signed($unsigned(reg523)));
              reg618 <= (^(~&$unsigned($signed($unsigned((7'h41))))));
              reg619 <= ((7'h4e) ^ (wire476[(1'h1):(1'h1)] ?
                  ($signed((+reg501)) ?
                      $unsigned($signed(wire483)) : (wire476[(4'hd):(4'hd)] == (reg547 ?
                          reg525 : wire478))) : (8'hbf)));
              reg620 <= reg595[(4'ha):(3'h6)];
            end
          else
            begin
              reg615 <= $unsigned(($signed(reg511[(4'h9):(1'h0)]) < $unsigned(wire564[(1'h1):(1'h1)])));
              reg616 <= $unsigned((^~wire485[(4'hb):(3'h6)]));
            end
          reg621 <= wire492[(4'hb):(3'h7)];
          reg622 <= reg515[(1'h1):(1'h0)];
          if ((~&$unsigned({reg594[(4'h8):(3'h6)]})))
            begin
              reg623 <= (reg504 ? (!(&{reg524[(5'h17):(4'ha)]})) : reg553);
              reg624 <= (reg595 ?
                  $signed($unsigned(reg500[(2'h3):(1'h1)])) : $signed(reg578));
              reg625 <= {($unsigned((8'hb4)) < reg527[(4'hf):(3'h7)]),
                  $signed((^{(reg538 ^ reg577)}))};
              reg626 <= ((^$unsigned((reg515 == (-reg547)))) ^ reg558[(4'hf):(2'h3)]);
            end
          else
            begin
              reg623 <= ({{reg497, reg542}} ?
                  ((($unsigned((7'h41)) ?
                          $signed(reg535) : reg522[(4'ha):(1'h0)]) + $unsigned($unsigned(reg538))) ?
                      reg592[(4'h8):(4'h8)] : ((8'ha2) ?
                          reg597 : ((reg527 & reg514) ?
                              $signed(wire485) : (8'ha5)))) : ($unsigned(({wire475,
                      (8'had)} < (reg589 && reg506))) || reg610[(5'h18):(3'h4)]));
              reg624 <= (&$unsigned(reg506));
              reg625 <= ({$signed($unsigned($unsigned(wire485))),
                      (+$signed($signed((8'hba))))} ?
                  (reg558 ? reg521 : (7'h48)) : reg501[(4'hd):(2'h2)]);
              reg626 <= $unsigned($signed((wire564[(2'h2):(1'h1)] < reg593[(1'h0):(1'h0)])));
            end
        end
    end
  assign wire627 = $unsigned(reg540[(1'h0):(1'h0)]);
  assign wire628 = wire484[(5'h14):(3'h7)];
  assign wire629 = (~&(^{(~^reg538[(1'h1):(1'h0)])}));
  assign wire630 = {{(|reg520)}, $unsigned(reg534[(1'h0):(1'h0)])};
  assign wire631 = ({reg583,
                       $unsigned(($unsigned(reg615) ?
                           (!reg502) : wire480[(3'h6):(2'h3)]))} << reg560[(1'h1):(1'h0)]);
  assign wire632 = {reg510[(1'h0):(1'h0)],
                       $unsigned($signed(((reg583 ~^ wire482) << reg499[(2'h2):(1'h0)])))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module199
#(parameter param469 = ((8'hb3) == ((-((~&(7'h42)) ? ((7'h49) ? (8'hbb) : (8'hbf)) : ((7'h43) >>> (8'ha2)))) ? (~|(+((8'hac) != (8'ha1)))) : ((((8'ha4) ? (8'hb0) : (8'hbf)) != ((7'h46) ? (7'h44) : (8'had))) ? ({(8'hb3)} ^ (|(8'hbc))) : ((|(8'hb9)) ? (+(8'hbb)) : ((8'ha6) <<< (8'h9e)))))), 
parameter param470 = (-(({(7'h44), (param469 >> param469)} < param469) || (param469 - (-(param469 ? param469 : param469))))))
(y, clk, wire203, wire202, wire201, wire200);
  output wire [(32'he6a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire203;
  input wire [(5'h15):(1'h0)] wire202;
  input wire signed [(4'hd):(1'h0)] wire201;
  input wire [(4'h8):(1'h0)] wire200;
  wire [(5'h19):(1'h0)] wire468;
  wire [(5'h14):(1'h0)] wire467;
  wire signed [(5'h14):(1'h0)] wire403;
  wire signed [(5'h1a):(1'h0)] wire402;
  wire [(5'h13):(1'h0)] wire401;
  wire [(5'h13):(1'h0)] wire400;
  wire signed [(5'h11):(1'h0)] wire399;
  wire signed [(4'h8):(1'h0)] wire398;
  wire signed [(3'h5):(1'h0)] wire351;
  wire signed [(2'h2):(1'h0)] wire294;
  wire signed [(2'h2):(1'h0)] wire293;
  wire [(3'h7):(1'h0)] wire292;
  wire signed [(3'h5):(1'h0)] wire291;
  wire [(4'ha):(1'h0)] wire290;
  wire signed [(5'h12):(1'h0)] wire289;
  wire signed [(4'hc):(1'h0)] wire288;
  wire [(5'h1a):(1'h0)] wire287;
  wire [(3'h4):(1'h0)] wire286;
  wire [(4'h9):(1'h0)] wire285;
  wire [(5'h13):(1'h0)] wire284;
  wire signed [(4'h8):(1'h0)] wire204;
  reg signed [(5'h13):(1'h0)] reg466 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg465 = (1'h0);
  reg [(3'h5):(1'h0)] reg464 = (1'h0);
  reg [(5'h19):(1'h0)] reg463 = (1'h0);
  reg [(4'hf):(1'h0)] reg462 = (1'h0);
  reg [(3'h6):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg459 = (1'h0);
  reg [(4'ha):(1'h0)] reg458 = (1'h0);
  reg [(3'h5):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg456 = (1'h0);
  reg [(4'hf):(1'h0)] reg455 = (1'h0);
  reg [(5'h10):(1'h0)] reg454 = (1'h0);
  reg [(5'h15):(1'h0)] reg453 = (1'h0);
  reg [(5'h11):(1'h0)] reg452 = (1'h0);
  reg [(5'h13):(1'h0)] reg451 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg450 = (1'h0);
  reg [(3'h4):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg448 = (1'h0);
  reg [(5'h19):(1'h0)] reg447 = (1'h0);
  reg [(4'ha):(1'h0)] reg446 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg445 = (1'h0);
  reg [(5'h16):(1'h0)] reg444 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg442 = (1'h0);
  reg [(5'h10):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg440 = (1'h0);
  reg [(5'h16):(1'h0)] reg439 = (1'h0);
  reg [(2'h2):(1'h0)] reg438 = (1'h0);
  reg [(5'h10):(1'h0)] reg437 = (1'h0);
  reg [(4'h9):(1'h0)] reg436 = (1'h0);
  reg [(4'h9):(1'h0)] reg435 = (1'h0);
  reg [(5'h18):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg432 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg431 = (1'h0);
  reg [(3'h7):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg429 = (1'h0);
  reg [(5'h14):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg426 = (1'h0);
  reg [(5'h10):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg423 = (1'h0);
  reg [(3'h5):(1'h0)] reg422 = (1'h0);
  reg [(5'h14):(1'h0)] reg421 = (1'h0);
  reg [(5'h12):(1'h0)] reg420 = (1'h0);
  reg [(4'he):(1'h0)] reg419 = (1'h0);
  reg [(4'he):(1'h0)] reg418 = (1'h0);
  reg [(4'hc):(1'h0)] reg417 = (1'h0);
  reg [(4'hb):(1'h0)] reg416 = (1'h0);
  reg [(3'h7):(1'h0)] reg415 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg413 = (1'h0);
  reg [(3'h4):(1'h0)] reg412 = (1'h0);
  reg [(5'h12):(1'h0)] reg411 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg410 = (1'h0);
  reg [(5'h19):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg407 = (1'h0);
  reg [(5'h15):(1'h0)] reg406 = (1'h0);
  reg signed [(4'he):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg404 = (1'h0);
  reg [(2'h3):(1'h0)] reg397 = (1'h0);
  reg [(3'h7):(1'h0)] reg396 = (1'h0);
  reg [(5'h19):(1'h0)] reg395 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg394 = (1'h0);
  reg [(5'h10):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg392 = (1'h0);
  reg [(3'h6):(1'h0)] reg391 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg390 = (1'h0);
  reg [(5'h17):(1'h0)] reg389 = (1'h0);
  reg [(5'h10):(1'h0)] reg388 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg387 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg386 = (1'h0);
  reg [(4'hd):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg384 = (1'h0);
  reg [(5'h14):(1'h0)] reg383 = (1'h0);
  reg [(5'h1a):(1'h0)] reg382 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg381 = (1'h0);
  reg [(5'h10):(1'h0)] reg380 = (1'h0);
  reg [(3'h4):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg378 = (1'h0);
  reg [(4'ha):(1'h0)] reg377 = (1'h0);
  reg [(3'h6):(1'h0)] reg376 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg375 = (1'h0);
  reg [(3'h5):(1'h0)] reg374 = (1'h0);
  reg signed [(4'he):(1'h0)] reg373 = (1'h0);
  reg [(4'he):(1'h0)] reg372 = (1'h0);
  reg [(5'h10):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg370 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg [(4'hd):(1'h0)] reg368 = (1'h0);
  reg [(4'h9):(1'h0)] reg367 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg365 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg364 = (1'h0);
  reg [(2'h3):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg361 = (1'h0);
  reg [(5'h14):(1'h0)] reg360 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg359 = (1'h0);
  reg [(2'h3):(1'h0)] reg358 = (1'h0);
  reg [(5'h16):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg356 = (1'h0);
  reg [(4'h9):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg [(2'h2):(1'h0)] reg350 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg348 = (1'h0);
  reg [(5'h16):(1'h0)] reg347 = (1'h0);
  reg [(3'h4):(1'h0)] reg346 = (1'h0);
  reg [(4'hc):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg344 = (1'h0);
  reg [(2'h3):(1'h0)] reg343 = (1'h0);
  reg [(5'h18):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg341 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg339 = (1'h0);
  reg [(5'h14):(1'h0)] reg338 = (1'h0);
  reg [(5'h11):(1'h0)] reg337 = (1'h0);
  reg [(4'hc):(1'h0)] reg336 = (1'h0);
  reg [(3'h5):(1'h0)] reg335 = (1'h0);
  reg signed [(4'he):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg333 = (1'h0);
  reg [(4'hd):(1'h0)] reg332 = (1'h0);
  reg [(4'hc):(1'h0)] reg331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg329 = (1'h0);
  reg [(5'h11):(1'h0)] reg328 = (1'h0);
  reg [(5'h13):(1'h0)] reg327 = (1'h0);
  reg [(3'h4):(1'h0)] reg326 = (1'h0);
  reg [(5'h15):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg323 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg321 = (1'h0);
  reg [(4'h8):(1'h0)] reg320 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg319 = (1'h0);
  reg [(5'h18):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg317 = (1'h0);
  reg [(4'hb):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg315 = (1'h0);
  reg [(3'h5):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg313 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg312 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg311 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg310 = (1'h0);
  reg [(2'h3):(1'h0)] reg309 = (1'h0);
  reg [(5'h18):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg306 = (1'h0);
  reg [(4'ha):(1'h0)] reg305 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg304 = (1'h0);
  reg signed [(4'he):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg302 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg301 = (1'h0);
  reg [(5'h16):(1'h0)] reg300 = (1'h0);
  reg [(4'he):(1'h0)] reg299 = (1'h0);
  reg signed [(4'he):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg297 = (1'h0);
  reg [(5'h1a):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg283 = (1'h0);
  reg [(4'hc):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg279 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg277 = (1'h0);
  reg [(5'h17):(1'h0)] reg276 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg275 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg274 = (1'h0);
  reg [(2'h2):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg271 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg270 = (1'h0);
  reg [(5'h10):(1'h0)] reg269 = (1'h0);
  reg [(5'h13):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg267 = (1'h0);
  reg [(3'h4):(1'h0)] reg266 = (1'h0);
  reg [(5'h1a):(1'h0)] reg265 = (1'h0);
  reg [(4'hc):(1'h0)] reg264 = (1'h0);
  reg [(4'he):(1'h0)] reg263 = (1'h0);
  reg [(4'hd):(1'h0)] reg262 = (1'h0);
  reg [(3'h7):(1'h0)] reg261 = (1'h0);
  reg [(5'h18):(1'h0)] reg260 = (1'h0);
  reg [(5'h10):(1'h0)] reg259 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg258 = (1'h0);
  reg [(5'h10):(1'h0)] reg257 = (1'h0);
  reg [(4'h9):(1'h0)] reg256 = (1'h0);
  reg [(4'hf):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg254 = (1'h0);
  reg [(4'hc):(1'h0)] reg253 = (1'h0);
  reg [(4'hf):(1'h0)] reg252 = (1'h0);
  reg [(5'h14):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg249 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg246 = (1'h0);
  reg [(2'h2):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg244 = (1'h0);
  reg [(5'h16):(1'h0)] reg243 = (1'h0);
  reg [(5'h14):(1'h0)] reg242 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg241 = (1'h0);
  reg [(5'h19):(1'h0)] reg240 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg239 = (1'h0);
  reg [(3'h4):(1'h0)] reg238 = (1'h0);
  reg [(5'h11):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg236 = (1'h0);
  reg [(3'h4):(1'h0)] reg235 = (1'h0);
  reg [(4'hc):(1'h0)] reg234 = (1'h0);
  reg [(4'h9):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg230 = (1'h0);
  reg [(3'h5):(1'h0)] reg229 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg228 = (1'h0);
  reg [(5'h18):(1'h0)] reg227 = (1'h0);
  reg [(4'he):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg225 = (1'h0);
  reg [(4'hf):(1'h0)] reg224 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg219 = (1'h0);
  reg [(3'h6):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg216 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg215 = (1'h0);
  reg [(5'h14):(1'h0)] reg214 = (1'h0);
  reg [(4'h9):(1'h0)] reg213 = (1'h0);
  reg [(4'hb):(1'h0)] reg212 = (1'h0);
  reg [(3'h6):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg208 = (1'h0);
  reg [(5'h10):(1'h0)] reg207 = (1'h0);
  reg [(4'h8):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg205 = (1'h0);
  assign y = {wire468,
                 wire467,
                 wire403,
                 wire402,
                 wire401,
                 wire400,
                 wire399,
                 wire398,
                 wire351,
                 wire294,
                 wire293,
                 wire292,
                 wire291,
                 wire290,
                 wire289,
                 wire288,
                 wire287,
                 wire286,
                 wire285,
                 wire284,
                 wire204,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 (1'h0)};
  assign wire204 = wire203[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      reg205 <= wire200[(3'h5):(3'h5)];
      if (wire201[(4'hd):(2'h2)])
        begin
          if ($signed(($signed(reg205) ?
              wire202 : {($signed(wire202) >= wire202)})))
            begin
              reg206 <= $unsigned((wire200[(3'h5):(1'h0)] ?
                  (^~$unsigned(wire202)) : (~^(((8'hb8) ? (8'ha3) : wire204) ?
                      (wire201 & wire202) : {wire200, wire204}))));
              reg207 <= {($signed($unsigned({wire203,
                      wire201})) ~^ $unsigned(reg205[(3'h7):(1'h0)])),
                  $signed(reg206[(3'h4):(2'h2)])};
              reg208 <= $signed(wire204[(1'h1):(1'h1)]);
              reg209 <= $signed((~|wire200[(3'h5):(3'h5)]));
              reg210 <= reg205[(5'h10):(4'hc)];
            end
          else
            begin
              reg206 <= (wire201[(3'h5):(1'h1)] ?
                  ((-(wire200[(2'h2):(2'h2)] ?
                          ((8'hbd) || wire200) : (~^wire203))) ?
                      reg209 : wire201) : (($unsigned($signed(reg210)) ?
                          $unsigned((~|wire202)) : $unsigned(wire201[(4'hc):(4'h9)])) ?
                      wire200[(2'h2):(2'h2)] : (^~((&wire203) <<< $signed(wire204)))));
            end
          if (reg210[(4'h8):(3'h7)])
            begin
              reg211 <= (((wire204[(3'h5):(2'h2)] ?
                          $signed($signed(reg208)) : wire200) ?
                      {(8'hb9)} : $unsigned($signed((^reg205)))) ?
                  (^~reg207) : wire200[(4'h8):(1'h1)]);
              reg212 <= $signed(reg209[(3'h5):(2'h2)]);
              reg213 <= $signed(wire202);
              reg214 <= reg205;
              reg215 <= ((reg213 == {(((7'h4a) + reg207) ?
                      $signed(reg210) : reg211[(2'h2):(2'h2)]),
                  {$signed(reg214),
                      reg213[(2'h2):(2'h2)]}}) <= reg208[(5'h11):(1'h0)]);
            end
          else
            begin
              reg211 <= (~$unsigned($signed($unsigned(reg214[(4'h9):(3'h4)]))));
              reg212 <= $signed({reg214});
            end
          if ((((~&reg214[(4'he):(2'h2)]) - (($signed((8'hb0)) <<< ((7'h45) ?
                  reg207 : (8'haa))) ?
              ($signed(reg214) ?
                  $unsigned(reg211) : (|wire201)) : ($unsigned(wire201) ?
                  (8'hbc) : $unsigned(reg215)))) != $unsigned($unsigned(wire200))))
            begin
              reg216 <= $signed(wire200[(2'h2):(1'h0)]);
              reg217 <= (7'h4e);
            end
          else
            begin
              reg216 <= $unsigned(wire202);
            end
          if ((~^{reg211}))
            begin
              reg218 <= $unsigned(((^~reg208[(2'h3):(1'h0)]) ?
                  reg206 : (reg210 * reg209)));
              reg219 <= $signed((~^(~(+reg207[(4'h8):(4'h8)]))));
              reg220 <= $signed($unsigned(reg216));
              reg221 <= (reg219[(1'h1):(1'h0)] <<< {$unsigned($signed($signed((7'h40)))),
                  {((reg215 ^ reg209) ^~ $unsigned(reg214))}});
              reg222 <= reg216;
              reg223 <= reg211;
            end
          else
            begin
              reg218 <= reg218;
              reg219 <= ((8'hac) ^~ $signed(wire202));
              reg220 <= wire201;
              reg221 <= reg212;
              reg222 <= ((wire202 == (-({(8'ha5)} ?
                  $unsigned(reg213) : (wire204 >>> (7'h4b))))) || $signed((((|wire204) ?
                      (8'hbb) : (reg209 ? (8'ha1) : (8'hb8))) ?
                  (^$signed((8'ha3))) : (!$signed((8'hb4))))));
            end
          reg224 <= $unsigned($signed($unsigned(reg219[(1'h1):(1'h0)])));
          reg225 <= (~|reg214[(4'h8):(1'h0)]);
        end
      else
        begin
          if ((~^(reg211[(1'h0):(1'h0)] + (7'h43))))
            begin
              reg206 <= reg214[(4'h8):(3'h7)];
            end
          else
            begin
              reg206 <= wire204;
              reg207 <= ((|reg206) && (((^(reg221 ?
                  reg210 : reg216)) | $signed((+reg219))) ^ reg214));
            end
        end
      if ((+wire200[(2'h3):(1'h0)]))
        begin
          reg226 <= $signed(($unsigned($unsigned(reg220)) ?
              (reg209[(4'ha):(2'h2)] >> ((~reg222) ?
                  (8'hae) : (reg207 ^~ reg211))) : ((7'h4e) < (~&(reg207 <= reg219)))));
          reg227 <= reg218[(3'h5):(2'h3)];
          if (((~$unsigned($unsigned((!reg223)))) ~^ wire202[(1'h1):(1'h1)]))
            begin
              reg228 <= {($unsigned((-$signed(reg223))) ?
                      ((reg205[(5'h11):(5'h11)] >= ((8'had) ?
                          (8'ha5) : reg224)) | (^(reg214 != wire202))) : (^wire201))};
              reg229 <= (~&(((7'h4c) ?
                  (^(reg214 << (8'ha2))) : $unsigned((~&(8'hae)))) >>> $signed(reg215)));
              reg230 <= ({(reg225[(5'h10):(4'hd)] ?
                          $unsigned(reg220) : $unsigned({wire204, (8'had)}))} ?
                  $signed($unsigned(($unsigned((8'ha8)) ^ reg222))) : ($signed({{reg217},
                      (reg206 <<< reg225)}) >= $unsigned($unsigned(reg209))));
              reg231 <= {reg208[(3'h6):(2'h2)]};
              reg232 <= $unsigned($signed($unsigned($unsigned((~reg207)))));
              reg233 <= ($unsigned((~|((reg230 * reg208) * (reg219 ?
                      reg212 : wire200)))) ?
                  ($unsigned(wire202) ?
                      (reg216[(3'h4):(1'h1)] ?
                          (+reg211) : wire203[(4'h9):(3'h7)]) : {$signed($unsigned(reg209)),
                          ($unsigned(reg206) ?
                              $signed(reg218) : reg223[(1'h1):(1'h1)])}) : reg209[(3'h4):(1'h0)]);
            end
          else
            begin
              reg228 <= ($unsigned(reg218[(2'h3):(2'h2)]) <= (reg227 ?
                  ({(reg216 == reg228)} ?
                      (~^$signed(reg205)) : $unsigned($signed(reg216))) : $signed(reg225[(3'h5):(2'h3)])));
              reg229 <= (~^(8'h9c));
              reg230 <= (8'ha0);
            end
          if ((~|(+reg207[(1'h0):(1'h0)])))
            begin
              reg234 <= ((((~&reg228) && {{(7'h45), reg205}}) ?
                      $signed(reg209[(5'h12):(4'hd)]) : reg232[(1'h1):(1'h0)]) ?
                  reg216 : $signed(((+$signed(reg210)) ~^ ($unsigned(reg223) << $signed(wire202)))));
              reg235 <= reg230[(4'h9):(3'h4)];
              reg236 <= reg228;
            end
          else
            begin
              reg234 <= ((&$signed($signed((reg217 == reg226)))) << $unsigned(((|wire200[(1'h1):(1'h1)]) ?
                  (8'hb3) : wire202)));
              reg235 <= $unsigned(((reg213[(1'h1):(1'h1)] <= (((7'h48) < reg221) ?
                      $signed(reg232) : reg222[(3'h5):(2'h2)])) ?
                  reg211 : $signed($signed($signed(wire204)))));
            end
          if (reg221)
            begin
              reg237 <= (((~reg221) << (((reg215 ~^ reg219) > $signed(reg232)) ?
                  (^~(~^reg210)) : wire204)) != ({(reg230[(4'hf):(1'h0)] || reg208),
                  wire202} ^~ reg220[(2'h2):(1'h0)]));
              reg238 <= ($signed(($unsigned(reg234) ?
                      ($unsigned(reg221) >= $signed(reg234)) : (|(reg233 ?
                          (8'haa) : reg226)))) ?
                  (reg234 ?
                      ($signed(reg229[(2'h3):(2'h2)]) ?
                          ((~|wire200) ?
                              (8'ha9) : reg235[(3'h4):(3'h4)]) : {reg229}) : (((reg231 >= reg221) ?
                              (8'hba) : reg219[(2'h2):(1'h0)]) ?
                          $unsigned({(7'h4a),
                              reg220}) : ((8'hb9) != (reg224 << (8'ha4))))) : $unsigned((!(reg217[(1'h1):(1'h1)] << (reg210 ^~ reg225)))));
              reg239 <= (|($unsigned(reg210) ?
                  (^$signed(wire200)) : ($signed((reg233 ? reg224 : reg221)) ?
                      $unsigned(reg237[(4'h9):(1'h0)]) : reg211)));
              reg240 <= reg223[(1'h0):(1'h0)];
              reg241 <= {$signed($signed($signed(reg226[(3'h7):(1'h1)]))),
                  ((-({reg234} ? reg215 : ((8'had) ? reg223 : reg207))) ?
                      ($signed($unsigned((8'ha2))) ?
                          (^(^reg206)) : reg228[(2'h3):(1'h1)]) : (($unsigned(reg232) ?
                              reg207 : reg228[(2'h3):(1'h0)]) ?
                          $signed(reg240[(4'hc):(1'h1)]) : reg227))};
              reg242 <= (reg235[(1'h1):(1'h1)] ?
                  (($signed(reg223) ?
                      $signed($unsigned((8'hbb))) : reg211) | (({reg213} + reg214) <<< {$unsigned(reg214)})) : $signed({{(~reg233),
                          $signed(reg226)},
                      $signed((reg219 == reg241))}));
            end
          else
            begin
              reg237 <= $signed((8'haf));
              reg238 <= reg240;
              reg239 <= (7'h48);
              reg240 <= (reg231 ?
                  reg217[(3'h5):(2'h3)] : (reg205 ?
                      $unsigned((!(^reg230))) : (8'ha1)));
            end
        end
      else
        begin
          if ((&(~|$signed($unsigned((reg206 > (7'h43)))))))
            begin
              reg226 <= $unsigned(($signed({$unsigned(reg211)}) ?
                  reg206 : (7'h4a)));
              reg227 <= (^reg207);
              reg228 <= (reg234 ? reg219 : wire201[(3'h4):(1'h1)]);
              reg229 <= (!wire200);
              reg230 <= reg228[(2'h3):(2'h2)];
            end
          else
            begin
              reg226 <= (^~reg241[(3'h4):(3'h4)]);
              reg227 <= (~^$signed((reg205[(4'he):(1'h0)] ~^ reg231[(2'h2):(1'h1)])));
              reg228 <= $unsigned(reg212);
              reg229 <= $unsigned($signed(reg222));
              reg230 <= $signed((^reg223));
              reg231 <= reg222;
            end
          reg232 <= {(reg230 && (reg210[(4'ha):(3'h7)] ?
                  (~|(wire200 >>> (8'hbf))) : {$unsigned(reg217),
                      $unsigned(reg219)}))};
        end
      if (reg215)
        begin
          if (reg239[(4'hb):(4'h8)])
            begin
              reg243 <= (reg241 ?
                  $signed((8'ha9)) : $unsigned(($signed((^~reg236)) ~^ (^~wire203[(3'h7):(3'h4)]))));
              reg244 <= (reg237 > $signed((reg214[(3'h4):(3'h4)] ?
                  {reg235[(3'h4):(1'h0)]} : {(~^(8'hbe)),
                      reg216[(4'h8):(1'h0)]})));
              reg245 <= reg229[(1'h0):(1'h0)];
              reg246 <= (7'h42);
              reg247 <= (&reg229[(3'h5):(3'h4)]);
            end
          else
            begin
              reg243 <= (({($unsigned(reg229) ? {reg243} : {reg229, reg225}),
                      $unsigned(reg235[(1'h1):(1'h0)])} ?
                  $unsigned($unsigned($unsigned(reg209))) : (^~{reg210})) << ((reg240[(4'hc):(4'hc)] && (reg242[(5'h11):(3'h7)] ?
                  {wire204,
                      reg221} : (reg242 <= (8'hbe)))) > reg214[(5'h14):(3'h6)]));
              reg244 <= (|reg212);
              reg245 <= reg217;
              reg246 <= {{$unsigned((-$signed((8'hb2))))}};
            end
        end
      else
        begin
          if (($signed({$signed((reg242 + (8'hb3)))}) >= reg212))
            begin
              reg243 <= ($unsigned((reg209[(1'h0):(1'h0)] >> (reg235 ?
                  {reg237, wire200} : (reg210 ?
                      reg224 : reg237)))) <<< $unsigned((((~&wire200) <= $signed(reg231)) ?
                  $signed(reg242[(4'he):(4'he)]) : reg233)));
            end
          else
            begin
              reg243 <= (!((wire204[(3'h4):(3'h4)] ?
                  (reg222 ?
                      reg209[(4'h9):(2'h3)] : $signed(reg220)) : reg231[(3'h6):(3'h6)]) ^ ((^reg238[(1'h0):(1'h0)]) ?
                  (&reg233) : reg229)));
              reg244 <= (!$signed(reg217));
              reg245 <= (reg219 <= $unsigned((reg213[(3'h6):(1'h0)] ?
                  {((7'h46) > reg240)} : reg223[(2'h2):(1'h0)])));
              reg246 <= ((~(reg222[(3'h4):(2'h3)] ?
                  (reg232 >>> reg215) : (reg207[(3'h7):(3'h5)] ^ (7'h45)))) & ($signed(($signed(wire201) ?
                      (reg206 << reg219) : (reg229 ? reg235 : reg245))) ?
                  $unsigned({{reg223}, $signed(reg238)}) : reg236));
              reg247 <= reg223[(1'h0):(1'h0)];
              reg248 <= (~&$signed(((|(!reg212)) + ((reg230 ^ reg240) && (reg216 ?
                  reg243 : reg212)))));
            end
          if (reg229)
            begin
              reg249 <= ($unsigned(reg247) ?
                  ($unsigned($unsigned($unsigned(reg229))) & reg209[(3'h7):(2'h3)]) : $unsigned(reg216));
              reg250 <= (!$signed((8'hbe)));
              reg251 <= $signed((+reg241[(4'h9):(4'h8)]));
              reg252 <= wire201[(4'hb):(4'hb)];
              reg253 <= {(reg209[(3'h7):(2'h3)] <= (reg244[(4'h9):(4'h9)] ?
                      (reg220 >> (8'ha2)) : (reg234[(4'h9):(3'h4)] < (^~reg222))))};
            end
          else
            begin
              reg249 <= $signed($unsigned(reg222));
              reg250 <= $signed(({$unsigned((|reg216)), reg235} ?
                  reg228 : {reg237[(3'h4):(2'h2)]}));
              reg251 <= $unsigned({{reg251}, reg253[(4'hc):(3'h7)]});
              reg252 <= $signed(reg235);
              reg253 <= $signed(reg233[(3'h7):(2'h3)]);
              reg254 <= (-reg234);
            end
          reg255 <= $signed($signed($signed((!reg245))));
          reg256 <= $unsigned(reg211);
          reg257 <= ($unsigned({reg218, {$signed((8'hb8))}}) ?
              {{$signed(reg208),
                      ((reg234 * reg243) ?
                          (reg232 ^ reg250) : (-reg214))}} : reg252[(3'h7):(1'h1)]);
          if ($signed(wire204[(1'h0):(1'h0)]))
            begin
              reg258 <= (~^(&(!{(reg212 & reg231),
                  (reg213 ? reg255 : reg232)})));
              reg259 <= reg243[(2'h2):(2'h2)];
              reg260 <= reg244;
              reg261 <= (^({((reg208 > reg216) ?
                          (reg218 >>> reg237) : $signed(reg217)),
                      reg221[(3'h6):(2'h3)]} ?
                  reg257[(4'hc):(4'hb)] : $signed($unsigned($unsigned(reg243)))));
              reg262 <= reg256[(2'h3):(2'h2)];
              reg263 <= ($unsigned((^~$unsigned(((8'h9d) ? reg214 : reg222)))) ?
                  $unsigned(($unsigned({(8'ha2),
                      reg256}) < (^~$unsigned(reg230)))) : reg208[(5'h10):(4'h9)]);
            end
          else
            begin
              reg258 <= ((8'ha4) ~^ (($unsigned($signed(reg217)) ^ {{(8'ha5),
                      wire201}}) && reg256));
              reg259 <= reg214;
              reg260 <= (wire201[(4'ha):(3'h6)] * ((reg208[(5'h11):(3'h5)] >> {(~^reg231)}) >= $signed($signed($unsigned(reg252)))));
              reg261 <= reg216[(4'hc):(3'h4)];
              reg262 <= reg206;
              reg263 <= {(+(((reg230 > reg212) ?
                      $signed(reg218) : (+reg254)) ^~ (~&$signed(reg258)))),
                  {(($unsigned(reg218) >>> $signed(reg227)) ?
                          reg240[(4'hf):(4'hf)] : reg208[(5'h10):(4'hf)]),
                      ($signed((reg234 ? reg222 : reg262)) ?
                          ((reg229 && reg243) ^ reg211) : ((~&(8'hb7)) == {reg263}))}};
            end
        end
      if ((($unsigned(((reg222 ?
          wire204 : reg222) & (reg253 || reg205))) <<< (~^((~^reg205) && {(7'h44),
          reg232}))) & (((^~$unsigned(wire200)) ?
              ((reg259 ^ reg241) ?
                  (reg213 == reg229) : ((7'h40) ?
                      reg260 : (8'hbb))) : wire203) ?
          $signed(reg259) : $unsigned(reg227[(4'hd):(4'ha)]))))
        begin
          if (reg251[(3'h4):(2'h2)])
            begin
              reg264 <= $unsigned($signed(reg208[(4'he):(3'h7)]));
              reg265 <= (~|reg210[(4'hf):(3'h5)]);
              reg266 <= (~|reg206[(3'h6):(2'h2)]);
              reg267 <= (^~$signed($signed($signed({reg239, reg220}))));
            end
          else
            begin
              reg264 <= $unsigned((reg208[(5'h12):(4'hf)] ?
                  {(reg260 ?
                          reg219[(1'h0):(1'h0)] : (reg218 ?
                              wire201 : reg237))} : reg230));
              reg265 <= reg258;
              reg266 <= (reg208 ? reg208 : {$signed(reg233)});
              reg267 <= wire202;
              reg268 <= reg217;
              reg269 <= (({reg206[(3'h5):(1'h0)],
                  ((+reg207) | {reg263})} < $unsigned(reg229)) >= {(~reg224[(4'hf):(3'h7)])});
            end
          reg270 <= $signed(reg236[(5'h12):(3'h4)]);
          if (reg247[(2'h3):(2'h3)])
            begin
              reg271 <= (~(($unsigned(reg246[(1'h1):(1'h0)]) * reg257[(4'hc):(1'h1)]) ?
                  reg258 : reg230));
              reg272 <= reg230[(4'h9):(4'h8)];
              reg273 <= (reg264 ?
                  reg223[(1'h1):(1'h1)] : {{$signed(reg219[(1'h1):(1'h0)]),
                          reg214[(4'hb):(2'h2)]}});
              reg274 <= (((((|(8'hae)) ?
                      reg255[(4'hb):(3'h6)] : $unsigned((8'ha6))) != reg247) ?
                  $unsigned({(|reg248), $signed(reg269)}) : ((8'hb9) ?
                      $unsigned({reg259}) : reg251)) ~^ reg208[(4'h8):(2'h3)]);
              reg275 <= reg235;
            end
          else
            begin
              reg271 <= ((reg216[(4'h9):(4'h9)] != (wire201 <= {$unsigned(reg226)})) ?
                  (reg269[(3'h5):(2'h2)] ?
                      $signed(($signed(reg256) ?
                          (wire201 ?
                              reg228 : reg265) : (~reg253))) : reg261[(3'h6):(1'h0)]) : reg216[(3'h4):(3'h4)]);
              reg272 <= (+(~^reg215));
            end
          reg276 <= reg253;
        end
      else
        begin
          if ((($unsigned((reg242[(4'hc):(3'h7)] <= $unsigned(reg232))) ?
                  $unsigned(reg252[(3'h6):(3'h6)]) : reg242[(4'h8):(3'h6)]) ?
              ($signed({(reg269 ? reg213 : reg218), wire202[(1'h1):(1'h0)]}) ?
                  {reg251[(4'ha):(1'h0)]} : $unsigned(reg237)) : $unsigned($unsigned(reg255[(4'hc):(2'h2)]))))
            begin
              reg264 <= reg239[(1'h0):(1'h0)];
              reg265 <= $signed(reg224);
              reg266 <= (($unsigned($signed($unsigned(reg270))) * (8'hb4)) ?
                  {($signed((reg250 & reg212)) ?
                          $unsigned(reg223[(2'h2):(1'h1)]) : ($signed(reg239) ^~ (+reg273))),
                      wire200[(1'h0):(1'h0)]} : $signed({(|{reg272, (8'hba)}),
                      ($unsigned(reg222) + reg274)}));
              reg267 <= {((-reg248[(4'hc):(2'h2)]) ?
                      (($signed(reg268) ~^ {(8'ha4)}) ?
                          (~&((7'h44) ? (8'ha6) : reg247)) : ((reg268 ?
                                  reg212 : reg224) ?
                              ((8'hac) >> reg224) : {reg271})) : $signed({(8'h9f),
                          reg236[(4'h8):(2'h2)]}))};
              reg268 <= reg234;
              reg269 <= wire201[(3'h6):(3'h6)];
            end
          else
            begin
              reg264 <= $signed(($signed(((reg259 + reg218) + reg223)) ?
                  (~$unsigned($unsigned(reg244))) : {(wire200[(2'h2):(1'h0)] ?
                          (|reg247) : (wire203 + (8'ha0)))}));
              reg265 <= reg212;
              reg266 <= $signed({({(reg244 >> (7'h41))} ?
                      {reg209[(3'h6):(1'h0)],
                          reg247} : $unsigned($unsigned(reg213)))});
              reg267 <= reg260;
              reg268 <= $signed((-$unsigned($unsigned(reg276[(3'h5):(2'h2)]))));
            end
          if ($signed(({$unsigned((reg219 > reg214))} ?
              (~|$signed((reg268 ? (8'hb2) : reg268))) : (&$unsigned((reg257 ?
                  reg221 : (7'h40)))))))
            begin
              reg270 <= (-$unsigned(((~|(reg224 ?
                  reg262 : reg219)) <= {$signed(reg238), $unsigned(reg270)})));
            end
          else
            begin
              reg270 <= $signed(reg260[(4'h9):(3'h5)]);
              reg271 <= $signed(reg213[(4'h8):(4'h8)]);
              reg272 <= $unsigned((8'hb6));
              reg273 <= $unsigned((((~|$signed(reg211)) ?
                  (reg266[(2'h3):(1'h0)] == $unsigned(reg271)) : reg241[(4'h8):(3'h7)]) || (~^wire201)));
              reg274 <= (reg216[(3'h6):(3'h4)] ?
                  reg207 : reg268[(4'he):(4'h9)]);
            end
          if (({(~|reg221)} ?
              reg274[(3'h4):(2'h3)] : (($signed((&wire200)) < $unsigned($unsigned(reg230))) | reg215)))
            begin
              reg275 <= (reg259[(2'h3):(2'h3)] ? reg214 : $unsigned((&reg256)));
              reg276 <= $unsigned({$signed(reg226)});
              reg277 <= reg248[(3'h4):(2'h2)];
              reg278 <= $unsigned(((+reg248[(1'h0):(1'h0)]) ?
                  reg234 : $unsigned((-$unsigned(reg270)))));
            end
          else
            begin
              reg275 <= ((~^((reg260 ?
                      $signed(reg210) : $signed((8'hbe))) | ((~&wire202) && ((8'h9e) >> reg274)))) ?
                  $unsigned(($unsigned(reg226) - ($signed(reg240) < $signed(reg275)))) : (reg215 + reg253[(3'h7):(1'h1)]));
              reg276 <= reg230[(1'h1):(1'h1)];
            end
          if (($signed((8'hb0)) - ((((reg246 ? reg215 : reg223) >>> ((8'had) ?
              reg252 : reg267)) + wire201) <= {((~|(8'hb1)) ?
                  (^reg243) : $unsigned(reg248)),
              ($signed(reg254) && reg272[(5'h11):(3'h6)])})))
            begin
              reg279 <= {(({reg237} == reg276[(5'h17):(1'h0)]) || reg264[(4'hb):(3'h4)]),
                  (((8'ha4) ?
                          $signed((|reg217)) : $signed((reg273 && reg270))) ?
                      reg249 : wire203[(4'h8):(4'h8)])};
              reg280 <= reg216[(3'h4):(1'h1)];
              reg281 <= reg237;
              reg282 <= $unsigned((reg274 ?
                  $unsigned((reg254[(5'h15):(5'h11)] ?
                      reg248[(2'h2):(2'h2)] : reg231[(3'h6):(1'h1)])) : ((^~$signed(reg260)) ?
                      $signed((reg267 <<< reg213)) : $signed({(8'hac)}))));
            end
          else
            begin
              reg279 <= $unsigned($unsigned((^((reg274 ?
                  reg278 : reg212) >= reg245[(1'h0):(1'h0)]))));
            end
          reg283 <= {(~^{{$signed(reg260), reg223[(2'h2):(2'h2)]},
                  ((-(8'ha9)) >> {reg245, reg244})}),
              ((~$signed((reg247 ? reg226 : reg208))) ?
                  (|(8'ha1)) : $signed(((^~reg256) ?
                      $signed(reg268) : (wire200 ? wire204 : reg233))))};
        end
    end
  assign wire284 = (!{{reg223, $signed((7'h44))}});
  assign wire285 = (+reg232);
  assign wire286 = (^reg228);
  assign wire287 = (!reg232);
  assign wire288 = (&(^$signed(reg260[(4'hf):(4'he)])));
  assign wire289 = (~($unsigned(reg242[(3'h6):(2'h3)]) ~^ $signed((((8'hac) | reg238) ?
                       $signed(reg251) : $unsigned((8'hba))))));
  assign wire290 = ((reg240 ?
                           $signed({(reg247 ? reg263 : reg281),
                               reg223[(1'h1):(1'h1)]}) : $signed({$unsigned(reg247),
                               reg252})) ?
                       (+$unsigned(reg276)) : ($unsigned(reg219[(2'h2):(1'h0)]) >= reg267));
  assign wire291 = (8'hb2);
  assign wire292 = {($signed($unsigned((-wire201))) ?
                           $unsigned($signed((wire203 && (7'h4d)))) : $signed(reg205))};
  assign wire293 = ($unsigned(reg226) ^~ reg228);
  assign wire294 = $signed(reg206[(3'h6):(3'h4)]);
  always
    @(posedge clk) begin
      reg295 <= $unsigned((($signed($unsigned(reg267)) ?
              $signed((wire293 ^~ reg225)) : (&(^~reg265))) ?
          (8'h9d) : reg265));
      if ((^reg241))
        begin
          if ({reg233[(3'h4):(3'h4)]})
            begin
              reg296 <= (^reg205);
            end
          else
            begin
              reg296 <= $signed(reg265[(4'hf):(1'h0)]);
              reg297 <= reg222;
              reg298 <= ((7'h4d) ?
                  (((&(reg281 ? (8'hb8) : reg273)) ?
                          (reg258 ?
                              $unsigned(wire292) : $unsigned(wire200)) : $signed(reg262[(4'hd):(3'h5)])) ?
                      ((((7'h44) ? reg222 : reg232) <= {reg238}) ?
                          ({(7'h49), reg276} ?
                              (~|reg240) : {reg282}) : reg280[(2'h2):(2'h2)]) : reg280) : wire204);
            end
        end
      else
        begin
          if ($signed(reg297[(4'hc):(3'h6)]))
            begin
              reg296 <= (wire289 + $unsigned($unsigned($unsigned((reg259 - (8'hbc))))));
            end
          else
            begin
              reg296 <= (~|(($signed(wire291[(2'h2):(1'h0)]) <= (~&$signed(reg225))) >> $signed(($signed((8'hb5)) >= {wire294}))));
              reg297 <= (&$unsigned((((wire284 ?
                  (8'haa) : wire291) * (wire287 >> reg244)) < reg263)));
              reg298 <= (($unsigned($signed((wire292 && reg230))) ?
                  (reg221 + $signed($signed(wire203))) : $unsigned(((reg258 ?
                          reg238 : reg279) ?
                      $signed(reg236) : reg274))) >>> wire201);
            end
          if (reg237)
            begin
              reg299 <= reg217;
              reg300 <= reg220;
              reg301 <= {({reg241[(1'h1):(1'h1)]} >= wire200[(3'h6):(1'h1)])};
              reg302 <= ($unsigned($unsigned((!(reg219 ?
                  reg213 : reg296)))) <<< (!$unsigned(reg283)));
              reg303 <= reg240;
              reg304 <= $unsigned(reg276[(2'h2):(1'h1)]);
            end
          else
            begin
              reg299 <= wire291;
              reg300 <= $unsigned($unsigned($signed((-reg255[(2'h2):(1'h0)]))));
              reg301 <= reg218;
              reg302 <= reg283;
              reg303 <= (~(~(8'hab)));
            end
          reg305 <= (^(((|$signed((8'ha5))) <<< (^$signed((7'h4c)))) - $unsigned(($unsigned(reg229) ?
              reg225 : $unsigned(reg279)))));
          reg306 <= $unsigned((reg229 || $signed(reg271)));
          if ((-reg295))
            begin
              reg307 <= reg303;
              reg308 <= $unsigned(($signed({reg275[(2'h2):(2'h2)]}) >= $signed(($signed(reg220) || $signed(reg240)))));
              reg309 <= ($unsigned({(~reg255),
                  ($signed(reg237) ?
                      $signed(reg223) : $signed(wire290))}) > ($signed(reg307) ?
                  $unsigned((~|(reg282 + reg216))) : (reg207[(4'hf):(2'h3)] < ($unsigned(reg252) != (reg267 != wire285)))));
              reg310 <= $signed((!$unsigned(((&reg208) ?
                  $signed((8'hb6)) : reg229))));
              reg311 <= $unsigned(reg278);
              reg312 <= $unsigned(reg268[(5'h13):(4'ha)]);
            end
          else
            begin
              reg307 <= (&(reg210[(2'h2):(2'h2)] && reg220[(2'h3):(1'h0)]));
              reg308 <= $signed(((~^(^~reg256[(3'h6):(3'h5)])) ?
                  reg271 : reg230));
              reg309 <= ({(($unsigned(reg268) ? (8'hbe) : reg264) ?
                          reg310 : reg252[(3'h6):(3'h5)])} ?
                  reg259[(4'he):(4'ha)] : (~|{reg222,
                      ((&reg299) | $unsigned(reg239))}));
            end
          reg313 <= (~(!{$signed((|reg281))}));
        end
      if ((~(8'hbd)))
        begin
          reg314 <= reg258;
          if (((^(-({wire285} ?
              ((7'h4d) ?
                  reg218 : (8'ha8)) : $unsigned(wire201)))) || $unsigned($signed(((reg278 <<< reg236) >>> (reg248 != (7'h47)))))))
            begin
              reg315 <= (reg238[(1'h0):(1'h0)] ?
                  reg300[(5'h13):(1'h1)] : (~^(8'had)));
              reg316 <= ((8'h9d) ^~ reg277[(5'h10):(3'h6)]);
            end
          else
            begin
              reg315 <= $signed($signed(reg272));
              reg316 <= $signed(reg222[(3'h6):(2'h3)]);
              reg317 <= reg269;
              reg318 <= $unsigned(reg301[(3'h6):(3'h4)]);
              reg319 <= reg265;
              reg320 <= (({((reg282 >= reg205) ? (7'h48) : (~&wire289)),
                          (wire204[(1'h1):(1'h1)] ?
                              (reg319 >> reg263) : (reg243 << reg224))} ?
                      $signed(((reg241 | wire285) ?
                          $unsigned(reg209) : (reg316 ^~ wire288))) : (($unsigned(reg234) ?
                          (reg279 ?
                              reg283 : reg240) : reg261[(3'h5):(3'h4)]) - (~reg211[(2'h2):(1'h0)]))) ?
                  ((reg229[(1'h0):(1'h0)] ?
                      reg297 : ($signed(reg244) ?
                          $unsigned(reg211) : ((8'ha5) << reg234))) >> (^~$signed($unsigned(reg312)))) : reg312[(1'h1):(1'h1)]);
            end
          if ($unsigned((8'hba)))
            begin
              reg321 <= $signed((|{(reg279 ? reg319[(2'h3):(1'h0)] : reg262),
                  $signed($signed(reg261))}));
              reg322 <= wire284;
              reg323 <= reg261[(1'h0):(1'h0)];
              reg324 <= (~(^~$unsigned($unsigned({reg279, reg281}))));
              reg325 <= reg256;
              reg326 <= (8'haf);
            end
          else
            begin
              reg321 <= ({(~(~$signed(wire286)))} || (reg253 || (((reg303 >= reg212) >= {reg228}) | reg245)));
              reg322 <= reg297;
            end
        end
      else
        begin
          if ((~|$signed((reg302 ?
              {(-(7'h47))} : (wire203 ?
                  (reg258 ? reg264 : reg226) : (~reg247))))))
            begin
              reg314 <= (8'ha2);
              reg315 <= $signed(reg208);
            end
          else
            begin
              reg314 <= ((({{(8'ha3), reg226}} * wire200[(3'h6):(1'h0)]) ?
                      $signed($signed(reg316)) : ((~&(-wire204)) ?
                          (~|reg280[(4'hd):(2'h3)]) : ((8'ha1) ?
                              (-reg279) : ((8'ha7) ? (8'hb1) : (8'hb8))))) ?
                  $signed($unsigned(((-wire293) >>> $unsigned((7'h4a))))) : reg321);
            end
          if ($unsigned($signed({$signed($signed((8'ha3)))})))
            begin
              reg316 <= $unsigned(reg236[(2'h3):(1'h1)]);
              reg317 <= (~|reg232[(2'h2):(1'h1)]);
              reg318 <= ((+(&$signed(reg315[(3'h4):(2'h2)]))) & ({reg306} ?
                  $unsigned(reg211[(1'h0):(1'h0)]) : reg314));
            end
          else
            begin
              reg316 <= $signed($signed(wire286));
              reg317 <= (~reg306[(2'h3):(2'h2)]);
              reg318 <= {reg306,
                  $signed((reg326 - $signed(reg313[(3'h4):(2'h3)])))};
              reg319 <= (|$signed($unsigned(({reg311, reg317} ^ (reg210 ?
                  reg212 : reg228)))));
              reg320 <= {(~|(((wire288 ? (8'haa) : reg283) ?
                      $unsigned(reg235) : $signed((7'h4e))) >= (reg256[(1'h1):(1'h0)] ?
                      reg207[(2'h3):(1'h0)] : $unsigned((7'h44)))))};
            end
          if ((reg265 < $unsigned((reg308[(3'h5):(2'h2)] ?
              ($unsigned(reg205) ?
                  (reg311 ?
                      reg226 : reg247) : ((8'hba) * reg299)) : reg283[(4'hc):(3'h6)]))))
            begin
              reg321 <= (-(^(|reg253[(1'h1):(1'h0)])));
              reg322 <= reg243[(1'h0):(1'h0)];
              reg323 <= reg239[(4'hd):(4'hc)];
            end
          else
            begin
              reg321 <= $signed($unsigned($signed($unsigned((~^reg251)))));
              reg322 <= ((reg312 + $signed({(~&reg247),
                  reg256})) > ((wire294[(2'h2):(1'h1)] ?
                      reg218[(3'h6):(1'h1)] : ({reg300} ?
                          ((7'h4d) ? reg265 : reg222) : $unsigned(reg326))) ?
                  (^~((reg248 ? (8'hb8) : wire284) << (reg233 ?
                      reg275 : (8'haf)))) : reg300[(4'hb):(4'hb)]));
              reg323 <= reg300;
              reg324 <= (($unsigned((^~$unsigned(reg325))) & $signed(({reg260,
                      reg299} ?
                  reg320[(1'h1):(1'h0)] : reg245))) & $unsigned(reg213[(4'h8):(3'h7)]));
              reg325 <= $unsigned(reg322);
              reg326 <= $signed($unsigned((~&(reg312[(2'h2):(1'h1)] ?
                  ((8'hb4) || wire284) : (reg314 ^ reg266)))));
            end
          reg327 <= reg300;
        end
      reg328 <= (~(7'h42));
      reg329 <= ((~&$signed(($unsigned((7'h45)) ?
          (reg210 >>> reg245) : (&reg225)))) ~^ {reg271[(3'h4):(2'h3)],
          $signed($signed($signed(reg249)))});
    end
  always
    @(posedge clk) begin
      reg330 <= {(!{$unsigned(reg261)}), (&reg303[(4'ha):(3'h4)])};
      reg331 <= $unsigned(reg268);
      reg332 <= $unsigned((8'ha0));
      reg333 <= $signed((~&reg258));
      if ((wire291 < $signed((~|{(reg277 ^~ reg271), reg276}))))
        begin
          if ((8'ha1))
            begin
              reg334 <= (!reg264[(1'h0):(1'h0)]);
              reg335 <= ((7'h4e) > ((-(|(~|reg239))) <= ((^(-(8'ha8))) ?
                  reg273[(2'h2):(1'h1)] : $unsigned((8'hb0)))));
              reg336 <= reg262;
              reg337 <= reg262[(2'h2):(2'h2)];
              reg338 <= $unsigned(wire284[(5'h12):(5'h11)]);
              reg339 <= {(&$unsigned(((wire204 + (7'h46)) ?
                      (~reg295) : $signed(reg338)))),
                  reg311[(4'h8):(3'h7)]};
            end
          else
            begin
              reg334 <= $unsigned(reg251);
              reg335 <= ((|$signed((!(^reg230)))) ?
                  $signed({($signed(reg236) ?
                          $unsigned(reg205) : (reg316 >> reg206))}) : (^~{(reg223 & $signed(reg323))}));
            end
          reg340 <= reg261;
          reg341 <= reg230[(3'h7):(1'h1)];
          reg342 <= {$unsigned((8'ha3))};
        end
      else
        begin
          if ($unsigned($unsigned($signed($signed({reg253})))))
            begin
              reg334 <= (reg276[(4'hf):(3'h5)] || ((((7'h4d) ?
                      reg216[(4'ha):(3'h4)] : reg262[(4'h8):(3'h6)]) ^ ({wire201} ?
                      wire294 : reg207)) ?
                  (reg296[(3'h6):(2'h2)] ?
                      $unsigned(reg205) : reg326[(2'h3):(2'h3)]) : {((|wire201) - reg257),
                      ($signed(reg257) | ((7'h42) && reg225))}));
              reg335 <= reg237;
            end
          else
            begin
              reg334 <= ((|$unsigned($unsigned($signed(reg227)))) ?
                  reg235[(1'h0):(1'h0)] : reg257[(2'h2):(1'h1)]);
              reg335 <= reg239[(1'h1):(1'h1)];
            end
          if ($signed(({$unsigned((reg266 == reg242))} > $unsigned(reg339))))
            begin
              reg336 <= ($unsigned(($unsigned($unsigned(wire291)) ?
                  (reg211[(1'h0):(1'h0)] ?
                      (reg250 ?
                          wire284 : reg240) : reg298[(2'h2):(2'h2)]) : $signed(wire288))) > {reg314[(3'h4):(3'h4)]});
              reg337 <= reg280;
              reg338 <= (8'hbe);
              reg339 <= $unsigned(($signed($unsigned((7'h4e))) == reg298[(3'h7):(1'h0)]));
              reg340 <= reg304;
              reg341 <= $signed($signed(reg317[(4'hc):(4'ha)]));
            end
          else
            begin
              reg336 <= reg306;
              reg337 <= $signed(($unsigned($signed(reg328[(4'hc):(4'hc)])) ?
                  (|$signed($signed((8'hb3)))) : {(^~(&reg262)),
                      (wire200 >> reg296)}));
              reg338 <= (wire285 ?
                  ((|((reg232 ? reg312 : reg208) ^ {reg295,
                      wire286})) <= reg340) : $unsigned($unsigned(($unsigned(reg304) | wire288))));
              reg339 <= {{((~^{reg211}) ?
                          $signed((~&reg238)) : (((8'ha3) ? reg315 : (8'ha6)) ?
                              (7'h4b) : reg269))},
                  reg237};
              reg340 <= ($signed((reg314 ?
                  ({reg331} ?
                      (reg326 ?
                          reg304 : reg211) : $signed((8'hb3))) : {(reg267 ?
                          reg300 : wire289),
                      $unsigned(wire203)})) ^ reg241);
            end
          if (((((reg305[(3'h7):(3'h4)] ?
                  $unsigned(reg279) : (&reg258)) * reg315) ?
              reg306[(1'h0):(1'h0)] : {$unsigned({wire288,
                      reg234})}) <= $unsigned({reg216[(1'h0):(1'h0)]})))
            begin
              reg342 <= $signed(reg276);
            end
          else
            begin
              reg342 <= ($unsigned($unsigned($unsigned((reg320 ?
                  wire285 : reg233)))) <= reg297);
              reg343 <= (&(7'h41));
              reg344 <= ((8'ha4) > (($unsigned((reg295 ? wire201 : wire289)) ?
                      (~&(reg279 + reg295)) : $unsigned($signed((8'hbc)))) ?
                  $signed(({reg298} ?
                      ((8'haa) ?
                          reg207 : reg279) : $signed(reg222))) : wire285[(2'h2):(2'h2)]));
              reg345 <= wire285;
            end
          if ((($unsigned((~$signed(reg245))) <<< ($signed($signed(reg308)) ?
                  ($signed(reg260) * (-wire293)) : reg297[(4'ha):(3'h6)])) ?
              $signed($unsigned($signed($signed((8'hac))))) : {reg345[(2'h3):(1'h0)],
                  reg230[(4'hd):(3'h5)]}))
            begin
              reg346 <= (reg244 ?
                  ($unsigned($unsigned((^~reg246))) ?
                      reg221[(3'h7):(3'h5)] : reg220[(2'h3):(1'h1)]) : reg240);
              reg347 <= reg300;
            end
          else
            begin
              reg346 <= reg255[(2'h3):(1'h1)];
              reg347 <= $unsigned(reg299[(1'h0):(1'h0)]);
              reg348 <= reg319;
              reg349 <= (reg239[(5'h10):(4'hb)] ?
                  ({{(8'hbf)},
                      $signed($signed(wire288))} <<< (~&((8'ha0) - reg332))) : (|({{reg245},
                      ((7'h4c) ? reg295 : reg277)} || reg216)));
              reg350 <= (reg226[(4'hb):(1'h0)] ?
                  ((8'hb8) ?
                      reg342[(5'h10):(3'h4)] : ({(~|reg318),
                          (^~(8'hb0))} | ((8'hbe) >> (reg266 | reg233)))) : (7'h4e));
            end
        end
    end
  assign wire351 = (!$unsigned(({reg317, {reg236}} ?
                       reg226[(4'hb):(3'h7)] : (|(wire292 >> reg283)))));
  always
    @(posedge clk) begin
      reg352 <= $signed($signed(wire286[(2'h2):(1'h1)]));
      if ($unsigned({$signed((reg223 ?
              $unsigned(reg223) : (reg308 ~^ (7'h46)))),
          $unsigned((~&$signed(reg346)))}))
        begin
          if (reg250)
            begin
              reg353 <= (+{$unsigned($signed($signed((8'hb9))))});
              reg354 <= ($unsigned((~((reg323 && reg212) ?
                  $signed(wire204) : (reg343 ? reg320 : reg270)))) || reg304);
              reg355 <= $signed(((({reg264,
                  reg246} | $signed(reg238)) >>> $signed((^reg206))) >= (~^(|reg223[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg353 <= $unsigned(reg298);
              reg354 <= $signed((((8'hba) ?
                  reg257[(1'h0):(1'h0)] : (reg268 ?
                      reg269 : (reg271 >= reg222))) >>> (reg250 >= reg221[(3'h4):(2'h2)])));
              reg355 <= reg327[(5'h13):(5'h11)];
              reg356 <= reg316[(1'h1):(1'h1)];
            end
          if ($unsigned(((&((reg238 ? reg242 : reg224) | (reg312 ^ reg330))) ?
              (!(^reg300[(3'h6):(1'h1)])) : reg319)))
            begin
              reg357 <= (!(~reg252[(3'h6):(2'h3)]));
            end
          else
            begin
              reg357 <= $signed(($signed(($unsigned(reg248) && $unsigned(reg243))) << ($unsigned((reg342 ^~ reg277)) != $unsigned($signed((8'ha1))))));
              reg358 <= $unsigned($signed(reg346[(2'h3):(1'h0)]));
              reg359 <= $signed((|$signed(($unsigned(wire204) >= $unsigned(reg251)))));
              reg360 <= reg352;
            end
          if (($unsigned(((~&$unsigned(reg341)) <<< $signed($unsigned(reg353)))) ?
              (((8'had) ?
                  wire200[(3'h7):(3'h6)] : $unsigned($unsigned(reg325))) * reg281) : $signed((((reg315 ?
                  reg278 : wire294) ^ (~^reg277)) ^ $unsigned((~reg230))))))
            begin
              reg361 <= (8'hae);
              reg362 <= ($unsigned({(-reg318[(1'h0):(1'h0)]), (7'h47)}) ?
                  {(~&reg325[(4'h9):(2'h2)])} : (reg336 + $signed((&(|(7'h49))))));
              reg363 <= reg217;
              reg364 <= reg362[(4'ha):(4'ha)];
            end
          else
            begin
              reg361 <= ((reg252[(1'h0):(1'h0)] ^ ((~|reg301) ?
                  ($unsigned(reg274) ?
                      (reg301 >>> reg324) : reg303[(3'h5):(1'h1)]) : $unsigned((~|reg249)))) == reg309);
              reg362 <= (({(reg364 << ((8'h9e) >= (7'h47))),
                          reg248[(2'h3):(1'h1)]} ?
                      $signed($signed({(8'hab)})) : {$unsigned((~&reg219)),
                          reg224[(4'ha):(1'h1)]}) ?
                  ($unsigned((|(&wire204))) >>> $signed((^((7'h49) < reg335)))) : $signed(($signed($signed(reg269)) ?
                      $signed(reg258[(2'h3):(2'h3)]) : {{reg316}})));
              reg363 <= $signed((8'ha1));
              reg364 <= $signed(reg300);
              reg365 <= $unsigned((&({{reg303}, (-reg270)} ?
                  ($signed(reg343) > (reg217 & reg220)) : $signed($signed(wire289)))));
              reg366 <= ((+reg323) ^ reg219);
            end
        end
      else
        begin
          reg353 <= (~reg228[(3'h6):(3'h5)]);
          reg354 <= {{(reg310[(1'h0):(1'h0)] ?
                      reg262[(1'h0):(1'h0)] : reg348)}};
          if ($signed(reg334))
            begin
              reg355 <= $unsigned((+reg331[(4'h8):(3'h4)]));
              reg356 <= reg346[(2'h3):(1'h0)];
              reg357 <= ($signed({$unsigned({(8'h9f), reg357})}) ?
                  ({(7'h44), {$unsigned(reg243)}} > {reg212,
                      ({reg283, reg231} ? reg353 : wire286)}) : (!reg328));
              reg358 <= (&reg356);
            end
          else
            begin
              reg355 <= (!reg340[(1'h1):(1'h1)]);
              reg356 <= (|$unsigned(wire289[(1'h0):(1'h0)]));
            end
          reg359 <= reg355;
          if ((+(reg295 == (^reg349[(3'h5):(1'h1)]))))
            begin
              reg360 <= reg210;
            end
          else
            begin
              reg360 <= (&((wire288 ?
                  (reg355[(3'h7):(3'h4)] == (~^(8'ha9))) : (^(reg341 ?
                      reg331 : reg302))) ~^ $signed(wire291[(1'h0):(1'h0)])));
              reg361 <= reg328[(4'hb):(1'h0)];
              reg362 <= reg345;
              reg363 <= (^$unsigned((^~{(reg263 ? reg303 : (8'hbd)),
                  (reg347 >>> reg360)})));
            end
        end
      if ($signed($unsigned(reg272)))
        begin
          if ($unsigned((reg208[(3'h7):(1'h1)] <= $unsigned(((reg271 >> reg229) ?
              (reg244 ? reg300 : reg342) : $unsigned(reg330))))))
            begin
              reg367 <= reg318[(3'h6):(1'h0)];
            end
          else
            begin
              reg367 <= (^(-$unsigned($unsigned($signed(reg278)))));
              reg368 <= ($signed(reg270[(1'h0):(1'h0)]) ?
                  ((&reg281) ?
                      $unsigned(($signed(reg334) ?
                          (~&reg229) : $signed((7'h4a)))) : wire200[(2'h3):(2'h2)]) : reg252);
              reg369 <= (reg336[(2'h2):(1'h1)] ?
                  ((8'ha5) ?
                      reg266 : (reg255[(4'hd):(3'h6)] ?
                          (((7'h4e) ^~ reg214) ?
                              reg257 : (~reg313)) : (+$signed(reg355)))) : (|reg229[(3'h5):(2'h3)]));
            end
          if ($unsigned(({{((8'hbd) ? reg222 : reg275),
                      reg272[(1'h1):(1'h0)]}} ?
              ((reg214 != (wire292 ?
                  (7'h47) : (8'h9e))) ~^ {(reg318 | reg223)}) : (|$unsigned($signed(reg308))))))
            begin
              reg370 <= ({$unsigned(((reg277 ? (8'ha2) : reg230) ?
                      reg237[(5'h11):(4'h8)] : (reg318 * (8'h9d))))} ^~ (reg227[(3'h7):(3'h7)] <<< $signed($unsigned((^reg367)))));
            end
          else
            begin
              reg370 <= $unsigned((&{$unsigned((~|reg349)),
                  wire285[(2'h2):(1'h1)]}));
              reg371 <= (($signed($signed((reg233 >>> reg223))) <= $signed((7'h45))) != {$unsigned(reg232[(1'h1):(1'h1)]),
                  (~^({reg332, reg318} || reg295[(5'h14):(4'ha)]))});
              reg372 <= reg340;
            end
        end
      else
        begin
          if ((reg343[(2'h2):(2'h2)] ?
              ($unsigned(reg260[(4'hc):(3'h4)]) <<< (~|reg205)) : ((reg270[(1'h0):(1'h0)] & ($signed(reg349) ^ wire203[(1'h0):(1'h0)])) ?
                  reg213[(3'h6):(3'h4)] : (-{(+reg305), {(8'haa), wire292}}))))
            begin
              reg367 <= reg259;
              reg368 <= $unsigned(reg370[(5'h13):(4'h8)]);
            end
          else
            begin
              reg367 <= reg370[(4'ha):(4'ha)];
              reg368 <= $unsigned((($signed((reg267 | wire289)) ?
                      (&$signed(wire203)) : reg271) ?
                  $unsigned($signed($unsigned(reg267))) : wire290[(3'h5):(2'h3)]));
            end
          reg369 <= $unsigned(wire200);
          if ($signed($signed($signed({{reg232, reg322}}))))
            begin
              reg370 <= $signed((-reg232[(2'h2):(1'h0)]));
              reg371 <= (+$signed((((reg341 <<< reg261) + reg271[(2'h3):(2'h3)]) ~^ (reg269[(3'h7):(2'h2)] >= (reg236 ?
                  reg283 : (8'hbf))))));
              reg372 <= reg215[(1'h0):(1'h0)];
              reg373 <= $unsigned((!$unsigned((reg212 ?
                  wire291[(2'h2):(1'h1)] : reg305[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg370 <= (reg338 ?
                  $unsigned(reg219[(1'h0):(1'h0)]) : $unsigned(reg226));
            end
        end
      if (($unsigned((reg275 ^~ ({reg216, (8'ha6)} ?
              (wire286 << reg258) : $signed((8'hae))))) ?
          wire203[(4'h9):(3'h6)] : $unsigned(reg236[(5'h11):(4'h8)])))
        begin
          reg374 <= reg342;
          if (($unsigned($signed(reg370)) ?
              $unsigned({$signed((reg365 ? (8'hb1) : wire201)),
                  reg232}) : ({reg251[(4'hb):(3'h5)]} - $signed((reg347 ?
                  reg212 : $unsigned(reg233))))))
            begin
              reg375 <= (reg333[(4'h9):(1'h1)] ?
                  $unsigned($signed((+reg252))) : reg271[(1'h0):(1'h0)]);
            end
          else
            begin
              reg375 <= (^({(~&(8'hb1))} == reg281));
              reg376 <= ((reg230 ? (^~reg278[(1'h0):(1'h0)]) : reg339) ?
                  reg264[(4'h8):(3'h5)] : (~&((reg358[(1'h1):(1'h0)] << {reg373}) >= (((8'hbd) - reg260) < (reg305 ?
                      reg362 : reg344)))));
              reg377 <= $unsigned($unsigned((reg295 ?
                  (&$signed((8'ha5))) : ($signed(reg324) ?
                      reg320[(3'h7):(1'h1)] : reg278[(1'h1):(1'h1)]))));
              reg378 <= $signed({(reg209[(5'h12):(4'h8)] ?
                      reg322[(3'h4):(2'h2)] : reg275)});
              reg379 <= ($unsigned({$signed((reg256 ? reg335 : (8'ha7)))}) ?
                  {reg344[(3'h4):(2'h3)],
                      (reg344 & ($signed(reg360) ?
                          reg368[(4'h8):(3'h7)] : $unsigned(reg370)))} : $signed((!((7'h49) ?
                      reg214 : $signed(reg272)))));
              reg380 <= ($signed({{$signed(reg260)}}) ?
                  $signed($unsigned((!reg275))) : $signed(reg341[(4'hf):(1'h0)]));
            end
        end
      else
        begin
          reg374 <= (+(+$signed($unsigned(wire201))));
          reg375 <= reg226[(1'h0):(1'h0)];
          if (({(((^~reg258) >= $signed(reg341)) ?
                      reg375 : (|$signed((8'ha3))))} ?
              ($unsigned((reg301[(1'h1):(1'h0)] ?
                      reg268[(2'h2):(1'h0)] : reg208)) ?
                  reg218[(3'h4):(2'h2)] : (reg313 ?
                      (!reg341) : {$unsigned(reg280),
                          (~reg257)})) : {(~(!(reg354 ? reg221 : wire284)))}))
            begin
              reg376 <= reg314[(1'h1):(1'h0)];
              reg377 <= (wire293 ^~ reg229[(3'h5):(2'h3)]);
              reg378 <= (7'h48);
              reg379 <= (reg257[(3'h7):(3'h5)] & ($signed(((reg361 ?
                  reg355 : (8'hb5)) && $signed((8'ha6)))) | (reg373[(2'h2):(1'h1)] ?
                  $unsigned($signed(reg345)) : reg273[(1'h1):(1'h1)])));
              reg380 <= $signed((8'ha0));
              reg381 <= $signed(wire288[(3'h5):(1'h1)]);
            end
          else
            begin
              reg376 <= $unsigned($unsigned($unsigned((~&reg213[(2'h3):(1'h1)]))));
              reg377 <= reg349;
              reg378 <= $unsigned((+$signed($signed((+reg374)))));
            end
        end
      if ((~^(reg248 & reg215)))
        begin
          if (reg276)
            begin
              reg382 <= (^$signed($unsigned((reg251[(4'h9):(1'h1)] && {reg380}))));
              reg383 <= ($signed(reg375[(1'h0):(1'h0)]) ^~ (~|(reg362[(5'h17):(5'h17)] ?
                  reg377 : ($signed(reg305) ?
                      reg266[(1'h0):(1'h0)] : (reg344 ? reg355 : reg312)))));
              reg384 <= reg315;
              reg385 <= (8'haf);
              reg386 <= $signed(({reg375} ?
                  (((reg236 ^ reg225) > $unsigned(reg313)) ?
                      ((~^reg266) <= (!reg208)) : reg343) : reg297[(1'h1):(1'h1)]));
              reg387 <= reg331;
            end
          else
            begin
              reg382 <= {(reg359 - $unsigned((reg346 ?
                      $unsigned(reg263) : (reg304 == reg223)))),
                  (reg302[(4'hc):(2'h2)] < $unsigned(reg275))};
              reg383 <= reg233;
              reg384 <= reg381;
              reg385 <= {$signed(reg208[(2'h2):(1'h0)])};
              reg386 <= reg315;
              reg387 <= (8'had);
            end
          if (($signed(reg255) - (&$unsigned(reg302))))
            begin
              reg388 <= $unsigned($unsigned(reg344[(3'h7):(2'h3)]));
              reg389 <= $signed(reg317[(2'h3):(1'h0)]);
              reg390 <= $unsigned($unsigned($signed((8'hbf))));
              reg391 <= {{reg215[(2'h3):(1'h1)]}, reg210};
            end
          else
            begin
              reg388 <= (reg245 != reg263);
              reg389 <= (reg297[(2'h2):(2'h2)] || (|($unsigned(wire292) ?
                  (7'h49) : $signed(wire293[(2'h2):(2'h2)]))));
              reg390 <= $signed(((({reg228, reg227} ?
                          ((7'h49) ^~ reg230) : (&reg298)) ?
                      $unsigned((reg328 ?
                          reg350 : reg316)) : $unsigned($unsigned(reg364))) ?
                  $unsigned((reg280[(4'hd):(4'h8)] ?
                      $unsigned(reg324) : (reg205 || reg364))) : (+$signed((~^reg205)))));
            end
          if (reg212[(1'h0):(1'h0)])
            begin
              reg392 <= ($signed(reg366) <= reg333);
              reg393 <= $unsigned(reg212[(1'h0):(1'h0)]);
              reg394 <= (((wire294 <= $signed(reg239[(4'h8):(3'h4)])) < (($unsigned(reg229) + $unsigned(reg262)) < ((reg385 - reg258) ?
                      (reg261 < wire294) : wire291[(1'h0):(1'h0)]))) ?
                  (($signed((reg252 != reg300)) ?
                      reg346[(1'h0):(1'h0)] : ((wire293 <= reg214) <<< (reg340 * reg365))) & (reg232 ?
                      $signed(wire285[(3'h7):(1'h0)]) : reg213[(4'h8):(2'h3)])) : (((-reg228[(4'h9):(2'h3)]) ?
                          (reg324[(4'he):(3'h7)] ?
                              (reg320 ?
                                  reg269 : reg217) : $unsigned((8'ha1))) : (reg233 ?
                              {reg309} : (reg367 << reg276))) ?
                      $unsigned($signed(reg337)) : $unsigned($signed({reg329,
                          reg390}))));
              reg395 <= (reg302[(1'h0):(1'h0)] ?
                  ($unsigned($unsigned(reg274[(4'hb):(4'hb)])) ?
                      $signed(reg272[(4'h9):(1'h1)]) : $signed($signed($signed(reg319)))) : reg367[(1'h0):(1'h0)]);
              reg396 <= (!(!$signed({reg319, reg231})));
            end
          else
            begin
              reg392 <= reg217;
              reg393 <= wire285[(4'h9):(3'h4)];
              reg394 <= reg217[(2'h3):(1'h0)];
              reg395 <= (+wire292);
              reg396 <= ($unsigned((!$signed((&reg377)))) >>> $unsigned($unsigned($signed({reg368}))));
            end
        end
      else
        begin
          if (reg355[(3'h6):(3'h4)])
            begin
              reg382 <= (8'ha9);
              reg383 <= (&($signed(((reg348 ? reg247 : reg253) ?
                      (reg276 ^~ wire293) : reg329[(3'h5):(2'h3)])) ?
                  ($unsigned($signed(reg342)) <= reg369) : {$unsigned(reg223[(2'h2):(1'h0)]),
                      (~^(~^reg385))}));
              reg384 <= {(reg248 ?
                      $signed({$unsigned(reg375),
                          $unsigned(reg323)}) : (((7'h4b) & reg319[(3'h4):(1'h0)]) <<< {(^~wire351)})),
                  reg206[(4'h8):(3'h7)]};
              reg385 <= $unsigned(reg384[(3'h4):(3'h4)]);
            end
          else
            begin
              reg382 <= $unsigned($signed((reg270 * reg232)));
              reg383 <= $unsigned($unsigned($signed(reg282[(3'h5):(2'h2)])));
              reg384 <= reg358;
              reg385 <= reg381;
            end
          reg386 <= ({$unsigned((+$unsigned((8'haf)))), reg207[(4'h8):(1'h0)]} ?
              (($unsigned(reg348) ?
                      $signed((-(7'h45))) : $unsigned({reg328, reg259})) ?
                  wire291 : reg264) : $signed((~|((reg389 ^~ reg316) ?
                  $unsigned(reg224) : (~^reg249)))));
          if ({$unsigned((8'h9f))})
            begin
              reg387 <= reg320[(4'h8):(4'h8)];
              reg388 <= $unsigned((reg394[(1'h1):(1'h1)] >= $unsigned((|{reg323}))));
              reg389 <= reg245[(1'h0):(1'h0)];
              reg390 <= (((($unsigned(reg344) || $unsigned(reg233)) ?
                  reg236 : (&{reg381})) >= ((!{wire201}) * wire293)) ^~ $signed({$unsigned(reg254),
                  ($signed(reg368) <<< $unsigned(reg223))}));
              reg391 <= reg367[(3'h5):(1'h0)];
              reg392 <= (reg214[(4'hf):(4'h8)] >>> (&reg270));
            end
          else
            begin
              reg387 <= (reg283[(4'hb):(2'h3)] >> {$unsigned((8'hb5)),
                  $unsigned(reg271)});
              reg388 <= reg382;
              reg389 <= ((8'h9d) | ($unsigned($signed((reg366 ?
                  (7'h4e) : reg350))) == (reg356[(4'h9):(2'h3)] ?
                  (reg386 >>> reg275[(3'h5):(3'h5)]) : {{reg368}})));
              reg390 <= ((^~($unsigned($signed(reg371)) >>> wire201[(4'h9):(1'h1)])) ^~ (reg206[(2'h3):(2'h2)] * $signed(reg326)));
              reg391 <= reg277[(1'h0):(1'h0)];
              reg392 <= reg263;
            end
          if ($signed(($signed(reg325[(3'h6):(3'h6)]) ?
              (^reg228) : {(~|(reg222 ? reg328 : reg264))})))
            begin
              reg393 <= (((reg301[(3'h4):(2'h2)] <= {reg384[(4'hb):(4'h9)],
                      (reg280 ?
                          reg250 : wire288)}) != $unsigned((!$unsigned(reg329)))) ?
                  ($signed($signed((~reg278))) ?
                      reg314 : {$unsigned(((8'hb6) ^ reg392))}) : $signed(reg226[(2'h3):(1'h0)]));
            end
          else
            begin
              reg393 <= (&reg396);
              reg394 <= (reg210[(5'h12):(3'h6)] != ((($unsigned(reg338) ?
                          (~|reg223) : wire293) ?
                      $unsigned(reg255) : $unsigned((~&reg205))) ?
                  {((-reg335) > (~^reg221)),
                      (reg362 ?
                          (7'h43) : (+reg243))} : $signed((~^(+reg382)))));
              reg395 <= $signed(wire290);
            end
        end
      reg397 <= $signed((~(reg278[(4'h9):(2'h2)] ?
          $signed($signed((7'h4a))) : (-((7'h4a) ? reg385 : (7'h4e))))));
    end
  assign wire398 = (reg393 | $signed($unsigned($unsigned((reg386 ?
                       wire284 : (8'had))))));
  assign wire399 = reg379[(1'h1):(1'h0)];
  assign wire400 = $signed({$unsigned(reg377), {reg309}});
  assign wire401 = (|reg225);
  assign wire402 = (^(wire399 ? reg367 : (~(^reg340))));
  assign wire403 = {{reg259[(4'hc):(1'h0)], reg311},
                       {reg345[(4'hc):(1'h0)], reg381[(5'h10):(1'h1)]}};
  always
    @(posedge clk) begin
      reg404 <= ((reg248[(4'h9):(1'h1)] ?
          reg211 : ((reg232[(1'h1):(1'h1)] ?
              $unsigned(reg328) : (reg392 < reg326)) << ((-reg308) ?
              wire286[(1'h1):(1'h1)] : reg299))) - $signed(reg269[(4'ha):(1'h0)]));
      if ((-(reg387[(1'h0):(1'h0)] ?
          (~reg233[(2'h3):(2'h2)]) : (wire291[(3'h4):(1'h0)] ?
              $signed($signed(wire291)) : $signed((reg327 ?
                  reg378 : reg374))))))
        begin
          if (reg370)
            begin
              reg405 <= $unsigned((~$unsigned(reg218[(1'h0):(1'h0)])));
              reg406 <= $signed(($unsigned((((8'haa) < reg212) ?
                      wire351[(1'h0):(1'h0)] : $unsigned(reg209))) ?
                  (&reg361[(3'h4):(2'h3)]) : $signed(($unsigned(reg324) ?
                      wire292[(3'h7):(1'h0)] : (reg254 ? reg304 : reg214)))));
              reg407 <= reg358;
              reg408 <= (reg338 | reg281);
              reg409 <= $signed($unsigned((+$unsigned((reg312 ?
                  reg313 : reg385)))));
              reg410 <= {(+reg297[(2'h3):(2'h3)]),
                  $signed($unsigned($signed(((8'hac) ? (7'h45) : reg396))))};
            end
          else
            begin
              reg405 <= ($signed(reg379[(3'h4):(1'h1)]) ?
                  ((|$unsigned((8'haf))) ~^ {((reg272 ?
                          wire288 : reg254) == (reg242 - reg279)),
                      $signed((reg377 >>> reg337))}) : $signed($unsigned($signed(reg377[(4'h9):(3'h7)]))));
              reg406 <= ($signed(reg281) || (^$signed(reg240)));
            end
          reg411 <= reg253[(3'h5):(3'h4)];
          if (($signed($unsigned((8'hba))) ?
              ((~reg359[(4'hc):(3'h7)]) <= ($unsigned($unsigned((8'h9c))) ?
                  $unsigned($signed((8'hb6))) : reg276[(2'h2):(1'h1)])) : ({($signed((8'h9e)) ?
                          reg271[(1'h1):(1'h1)] : (reg205 ? reg377 : reg349))} ?
                  (reg215[(2'h3):(1'h0)] ?
                      (reg319 == reg257[(3'h6):(3'h6)]) : $signed((reg255 > reg396))) : $signed(reg356))))
            begin
              reg412 <= ($signed($signed(((-reg262) ?
                      reg357[(5'h11):(4'hb)] : reg334[(4'h8):(1'h0)]))) ?
                  $unsigned(((reg260 ? (+reg259) : (-reg320)) ?
                      ((reg388 ? reg331 : reg257) ?
                          $unsigned(reg222) : ((7'h4d) ?
                              reg348 : wire284)) : $unsigned($unsigned(reg245)))) : (reg361[(3'h4):(3'h4)] ?
                      (reg320[(2'h2):(1'h0)] ?
                          (~(&reg331)) : (^(|reg348))) : $unsigned((!$unsigned(reg359)))));
              reg413 <= $unsigned((8'haa));
            end
          else
            begin
              reg412 <= ((~(($signed(reg374) >> {reg376,
                      reg329}) ^~ reg409[(5'h18):(3'h4)])) ?
                  reg253[(3'h5):(3'h4)] : (~&(+wire401)));
              reg413 <= $unsigned((((^~$signed(reg267)) + reg405[(3'h5):(1'h0)]) == reg394));
            end
        end
      else
        begin
          reg405 <= $unsigned($unsigned((((reg326 <= reg371) ?
              {reg321} : $signed(reg220)) >= (~&(&reg307)))));
        end
      if (($signed((reg302[(4'hd):(1'h1)] ?
          $signed(reg222[(4'hb):(1'h1)]) : wire202)) != (8'ha8)))
        begin
          reg414 <= reg320;
          if ({((((-(7'h47)) | (reg280 <<< reg348)) ?
                  $signed(reg267[(4'ha):(2'h3)]) : reg307) >>> (+((reg225 == reg363) ~^ wire289[(4'hf):(1'h1)])))})
            begin
              reg415 <= $unsigned($signed($unsigned($signed((reg245 == reg349)))));
            end
          else
            begin
              reg415 <= reg325;
              reg416 <= reg362[(5'h12):(5'h11)];
              reg417 <= (reg328 ?
                  ((reg340 >> $unsigned((+reg299))) < {$signed(reg223),
                      $signed((reg404 ? reg321 : reg235))}) : ((reg222 ?
                      reg236[(3'h7):(3'h6)] : reg216[(1'h1):(1'h0)]) <<< ((8'ha1) ?
                      $unsigned($unsigned(reg350)) : $unsigned(reg300[(5'h15):(4'h9)]))));
              reg418 <= (!reg332);
              reg419 <= (reg208 >>> $signed((^~($unsigned(reg395) ?
                  {reg386} : $signed(reg371)))));
              reg420 <= $unsigned((&wire398));
            end
          reg421 <= ((+reg247) ?
              $signed((^$signed(reg300))) : ($signed(reg263) - $signed(reg252)));
          reg422 <= ($unsigned((~wire200[(3'h4):(1'h1)])) < reg217);
          reg423 <= $signed({$signed(reg349)});
          if ((($unsigned((|$unsigned(reg414))) + reg346) ?
              (8'hbb) : $signed(($unsigned((^~reg237)) >> wire204[(2'h2):(1'h0)]))))
            begin
              reg424 <= (reg343 < (((!$signed(wire293)) ?
                  (~$signed(reg361)) : reg332[(4'hd):(4'hb)]) == reg271));
              reg425 <= {$signed($unsigned((7'h4b)))};
              reg426 <= ((~^$unsigned(({reg418, reg377} ?
                      $signed(reg376) : {reg421, reg419}))) ?
                  {(!$unsigned((-(8'hba))))} : reg315);
            end
          else
            begin
              reg424 <= ((reg312[(2'h2):(2'h2)] >= {($unsigned(reg230) < (8'hac))}) ?
                  $unsigned($unsigned((~|((7'h40) * (7'h4d))))) : reg361[(3'h4):(1'h0)]);
              reg425 <= reg326[(2'h2):(2'h2)];
              reg426 <= (~^{(+(^~reg337)), reg324[(4'hb):(3'h5)]});
              reg427 <= (~^$signed($unsigned(reg232)));
            end
        end
      else
        begin
          reg414 <= $unsigned((^(($unsigned((8'had)) >= wire398) ?
              ($unsigned(reg373) >> {reg421,
                  reg392}) : ((~^reg382) && reg212[(3'h6):(2'h2)]))));
          reg415 <= $signed((~^reg424));
          if ($unsigned($signed($unsigned(((reg325 ? reg384 : reg227) ?
              reg314 : reg276)))))
            begin
              reg416 <= reg425[(4'he):(4'hc)];
              reg417 <= $signed(reg313[(5'h19):(3'h5)]);
              reg418 <= reg331[(4'h8):(4'h8)];
              reg419 <= reg224;
            end
          else
            begin
              reg416 <= (8'hb4);
              reg417 <= (~^reg396[(2'h3):(2'h2)]);
              reg418 <= reg320[(2'h3):(2'h2)];
              reg419 <= $unsigned(($unsigned(($signed(reg312) ?
                      reg418 : (reg397 == (8'ha6)))) ?
                  reg334[(3'h4):(2'h2)] : (~&{(+reg240)})));
            end
          if ($unsigned($signed((reg394[(2'h2):(1'h0)] <<< reg238))))
            begin
              reg420 <= $signed((reg376[(2'h3):(1'h1)] >>> (&$signed((reg300 ?
                  (7'h44) : wire288)))));
            end
          else
            begin
              reg420 <= $unsigned((^~(reg264[(3'h7):(1'h1)] + ($unsigned(reg271) ?
                  reg348[(2'h3):(1'h1)] : $unsigned(reg382)))));
              reg421 <= ($signed(reg265[(3'h7):(3'h6)]) ^~ $unsigned((~$signed($signed(reg222)))));
              reg422 <= reg373[(3'h7):(2'h3)];
              reg423 <= reg242;
              reg424 <= (reg220[(2'h2):(1'h0)] ?
                  reg424[(5'h18):(4'ha)] : $unsigned((reg323 ?
                      (reg219[(1'h0):(1'h0)] ?
                          reg232 : ((8'hac) > reg247)) : (~^$unsigned(reg404)))));
              reg425 <= $signed(reg319[(1'h1):(1'h1)]);
            end
          reg426 <= $unsigned((&reg247));
        end
      reg428 <= (^($signed(reg388[(4'hf):(4'hb)]) ?
          (^reg323[(5'h13):(5'h11)]) : {$unsigned($signed(reg232)), reg337}));
      if (((reg325[(3'h6):(1'h0)] ?
          {($signed(reg207) ?
                  {reg324, (8'hb6)} : (wire201 ?
                      reg249 : (8'hb7)))} : $signed((7'h4a))) == reg257[(1'h1):(1'h0)]))
        begin
          reg429 <= reg356[(3'h6):(1'h1)];
          reg430 <= $signed($signed(({reg383[(4'hb):(3'h7)],
                  $unsigned(reg213)} ?
              (~|(8'hb7)) : (reg376 & (reg233 ? reg225 : reg345)))));
          if (((~|($unsigned(reg281[(4'hc):(3'h5)]) >> wire293)) < (reg219[(1'h1):(1'h1)] ?
              $signed($signed($signed(wire288))) : reg269)))
            begin
              reg431 <= (reg313 << reg244[(3'h6):(1'h0)]);
            end
          else
            begin
              reg431 <= ($signed({($signed((8'hb6)) ^~ (reg255 ~^ reg334)),
                      $signed($signed(reg338))}) ?
                  ($unsigned({((8'hb5) ? reg412 : wire288)}) ?
                      wire286[(1'h0):(1'h0)] : (((wire400 ?
                              reg378 : reg348) ~^ wire289) ?
                          (^~$unsigned(reg249)) : ((reg270 | reg348) || $unsigned(reg340)))) : (reg271[(2'h2):(1'h0)] ?
                      (+(-$unsigned(reg215))) : $signed(reg406[(3'h6):(3'h6)])));
              reg432 <= ((|reg239[(2'h3):(2'h3)]) < $unsigned(((~&$signed(reg246)) ?
                  (!reg273) : $unsigned({reg346, (8'hb2)}))));
              reg433 <= $signed($unsigned($unsigned((~reg396))));
            end
          reg434 <= ($signed({$unsigned($signed(wire398)),
                  (~|$unsigned((8'hac)))}) ?
              {(reg226 ?
                      (~&(wire351 ? (8'hab) : reg211)) : ($signed(reg425) ?
                          wire203[(4'hc):(4'h9)] : (^~(8'haf))))} : $unsigned(reg250[(2'h3):(2'h3)]));
          if (((!reg308) | (7'h44)))
            begin
              reg435 <= $signed(reg312);
              reg436 <= reg412[(2'h3):(2'h3)];
              reg437 <= {($signed(reg361) < $unsigned((8'haa)))};
              reg438 <= (reg427 * (((^~reg320[(3'h4):(1'h1)]) != ((-wire291) - reg257[(3'h5):(1'h0)])) ^ (8'h9c)));
              reg439 <= (^$unsigned($signed((reg345 << (wire204 * wire293)))));
            end
          else
            begin
              reg435 <= reg213;
              reg436 <= (~(8'hb6));
              reg437 <= $signed($signed($unsigned({(+(7'h42))})));
              reg438 <= ($unsigned($signed(({reg353,
                      reg381} + $unsigned(reg409)))) ?
                  reg212[(1'h0):(1'h0)] : reg218[(3'h6):(1'h1)]);
              reg439 <= reg302;
              reg440 <= $signed((~reg377[(3'h7):(3'h5)]));
            end
        end
      else
        begin
          if ((wire400 > ($unsigned(reg350) ?
              $unsigned($unsigned((reg335 == reg349))) : $signed((^~{wire288})))))
            begin
              reg429 <= ($unsigned(wire287[(4'hd):(1'h0)]) ?
                  (8'hb0) : $unsigned(reg356));
              reg430 <= (&$unsigned($unsigned($signed((!reg277)))));
              reg431 <= (+reg390[(3'h5):(1'h0)]);
            end
          else
            begin
              reg429 <= wire401;
            end
        end
      reg441 <= (|$unsigned(((^~$signed(reg276)) > reg315[(1'h1):(1'h0)])));
    end
  always
    @(posedge clk) begin
      if ($signed((~reg374[(3'h4):(1'h1)])))
        begin
          reg442 <= (($unsigned(reg430[(3'h7):(1'h1)]) | $signed({(-reg231)})) <<< (|reg354[(3'h4):(3'h4)]));
          reg443 <= ((($signed(wire293[(1'h0):(1'h0)]) ?
                  $unsigned(reg211[(1'h1):(1'h0)]) : (((8'hbc) ?
                      reg262 : reg380) > $signed(reg397))) ?
              reg240[(4'hc):(4'h8)] : $signed(((-(7'h4d)) ~^ ((8'hb9) ?
                  reg406 : reg427)))) <= (|(-($signed((7'h4a)) ?
              (reg297 ? reg392 : reg428) : (reg255 ? (7'h41) : reg268)))));
        end
      else
        begin
          reg442 <= (|$signed(reg312[(1'h0):(1'h0)]));
        end
      if (($unsigned({($signed((8'h9e)) << $signed(reg314)),
          ((reg261 ?
              reg225 : (7'h45)) && reg373[(4'he):(3'h7)])}) + reg240[(1'h1):(1'h0)]))
        begin
          reg444 <= reg231[(4'h9):(2'h3)];
          reg445 <= $unsigned({{((&reg329) ^~ (^reg419))}});
          if (reg396[(3'h6):(3'h4)])
            begin
              reg446 <= (~^$signed((-({reg358,
                  (8'hb7)} + (reg226 ~^ reg238)))));
              reg447 <= reg385[(4'hb):(4'h9)];
              reg448 <= reg257;
              reg449 <= (-(+$unsigned($unsigned((reg438 ? reg419 : wire200)))));
              reg450 <= {(~^reg252), $signed(reg329)};
              reg451 <= (reg364 <= (^wire398));
            end
          else
            begin
              reg446 <= (reg360 ?
                  (reg335 >> (reg314 ?
                      $signed($unsigned(wire201)) : $signed((|wire293)))) : reg251[(3'h7):(2'h3)]);
            end
          reg452 <= reg412;
          if (reg310[(2'h3):(2'h2)])
            begin
              reg453 <= (+((~$unsigned(((8'h9f) != reg389))) ?
                  (&reg411[(5'h10):(3'h6)]) : reg305[(2'h2):(1'h0)]));
              reg454 <= $unsigned((~reg312[(1'h1):(1'h1)]));
              reg455 <= ($unsigned(((reg244[(1'h0):(1'h0)] ?
                      $signed(reg261) : $signed(reg432)) | ($signed(reg215) < $signed(reg254)))) ?
                  $unsigned((~&$unsigned($signed(reg309)))) : (-$unsigned($signed(reg256))));
              reg456 <= ($signed({{(reg237 ? reg271 : reg231)},
                  $signed($unsigned((8'h9e)))}) < (((reg237 ?
                      $unsigned(reg409) : reg335[(1'h0):(1'h0)]) & (^(reg365 - reg222))) ?
                  ((reg305 ? (reg423 < (7'h4c)) : (reg370 ? reg342 : (7'h48))) ?
                      ((^~reg335) ?
                          reg434[(4'h8):(4'h8)] : (reg443 > (7'h4a))) : (|(-(8'hb6)))) : reg272));
              reg457 <= (~|$signed(reg415[(3'h4):(2'h3)]));
            end
          else
            begin
              reg453 <= ((&((|reg264[(1'h1):(1'h1)]) ?
                      reg362 : reg454[(3'h7):(3'h7)])) ?
                  reg438 : ((($unsigned((7'h4c)) ?
                          ((8'hb7) ?
                              wire292 : (8'hae)) : $signed(reg412)) && reg254) ?
                      reg364 : (((reg300 >= reg392) == (reg414 ?
                              reg305 : (8'hbb))) ?
                          $unsigned($signed(reg428)) : (reg377 ?
                              reg302[(3'h5):(1'h0)] : $signed(reg335)))));
            end
          if ($unsigned(reg339[(1'h1):(1'h1)]))
            begin
              reg458 <= reg279;
              reg459 <= ((-reg408[(3'h6):(3'h5)]) ?
                  (reg433 < reg235[(2'h3):(2'h2)]) : ({((^~reg358) && $unsigned(wire293)),
                      reg267[(4'ha):(3'h4)]} >> ($unsigned($unsigned(reg248)) * reg391)));
              reg460 <= reg322[(2'h2):(2'h2)];
              reg461 <= reg323;
              reg462 <= reg301;
              reg463 <= $signed(reg238[(1'h0):(1'h0)]);
            end
          else
            begin
              reg458 <= ($unsigned((reg411 ?
                  (reg303[(3'h7):(3'h7)] ?
                      (^~reg393) : (&reg228)) : reg355)) - reg450);
              reg459 <= (7'h46);
            end
        end
      else
        begin
          reg444 <= $unsigned(reg387[(3'h4):(2'h3)]);
        end
      reg464 <= ((reg270[(1'h0):(1'h0)] ?
          (reg240 ^~ reg274) : $signed(((reg259 == reg352) - $signed(reg383)))) <= (~reg336));
      reg465 <= (reg454[(1'h1):(1'h0)] ?
          $unsigned(reg433[(1'h1):(1'h0)]) : $unsigned(((~|reg305[(2'h2):(2'h2)]) ?
              $unsigned($unsigned(reg447)) : reg416)));
      reg466 <= ($unsigned($unsigned({(|reg210)})) ?
          reg392[(2'h2):(2'h2)] : (~|$signed($signed($signed(reg409)))));
    end
  assign wire467 = reg405;
  assign wire468 = $signed((wire399[(4'hb):(1'h1)] < reg452));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module187  (y, clk, wire192, wire191, wire190, wire189, wire188);
  output wire [(32'h21):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire192;
  input wire signed [(4'hc):(1'h0)] wire191;
  input wire [(5'h19):(1'h0)] wire190;
  input wire [(2'h3):(1'h0)] wire189;
  input wire signed [(4'hc):(1'h0)] wire188;
  wire signed [(3'h6):(1'h0)] wire196;
  wire signed [(3'h4):(1'h0)] wire195;
  wire signed [(3'h4):(1'h0)] wire194;
  wire [(5'h12):(1'h0)] wire193;
  assign y = {wire196, wire195, wire194, wire193, (1'h0)};
  assign wire193 = (((~|$signed((7'h44))) ?
                       ((~&wire188) ?
                           $unsigned({wire192}) : $unsigned((8'hb3))) : $unsigned(wire189[(2'h3):(2'h2)])) & (wire192 ?
                       (wire191[(2'h2):(1'h1)] ^~ wire192) : ($unsigned($signed(wire190)) >> (+wire192[(4'h9):(2'h3)]))));
  assign wire194 = ((($signed((|wire188)) ?
                               $signed(wire191[(3'h5):(1'h0)]) : $signed(wire192)) ?
                           $unsigned((~&(wire189 - wire189))) : (!(wire190 ^ (wire190 ?
                               wire193 : (8'hae))))) ?
                       $unsigned($signed($unsigned((wire190 | (7'h4e))))) : {$signed(wire191[(4'hc):(2'h2)])});
  assign wire195 = wire188;
  assign wire196 = wire195[(1'h1):(1'h1)];
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param997 = (&((&((~|(8'h9e)) ? (|(8'ha9)) : (~|(8'hba)))) ^ {(~((8'hb2) ? (8'h9e) : (8'ha4))), {{(7'h40), (8'ha4)}, (^~(8'h9c))}}))
, parameter param998 = param997 )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h63d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire0;
  input wire [(4'hf):(1'h0)] wire1;
  input wire [(4'he):(1'h0)] wire2;
  input wire signed [(2'h3):(1'h0)] wire3;
  input wire signed [(4'ha):(1'h0)] wire4;
  wire [(4'h9):(1'h0)] wire996;
  reg [(4'he):(1'h0)] reg995 = (1'h0);
  reg [(4'hd):(1'h0)] forvar994 = (1'h0);
  reg [(5'h15):(1'h0)] reg993 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg986 = (1'h0);
  reg [(5'h11):(1'h0)] forvar984 = (1'h0);
  reg signed [(4'he):(1'h0)] reg992 = (1'h0);
  reg [(4'hc):(1'h0)] reg991 = (1'h0);
  reg [(3'h5):(1'h0)] reg990 = (1'h0);
  reg [(5'h14):(1'h0)] reg989 = (1'h0);
  reg [(4'h8):(1'h0)] reg988 = (1'h0);
  reg [(4'hc):(1'h0)] reg987 = (1'h0);
  reg [(4'he):(1'h0)] forvar986 = (1'h0);
  reg [(4'hc):(1'h0)] reg985 = (1'h0);
  reg [(4'ha):(1'h0)] reg984 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg983 = (1'h0);
  reg [(5'h11):(1'h0)] reg982 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg980 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg979 = (1'h0);
  reg [(3'h5):(1'h0)] forvar978 = (1'h0);
  reg [(3'h6):(1'h0)] reg977 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar976 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg975 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg973 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg972 = (1'h0);
  reg [(5'h12):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg970 = (1'h0);
  reg [(3'h7):(1'h0)] forvar969 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar968 = (1'h0);
  reg [(4'hb):(1'h0)] reg967 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar966 = (1'h0);
  reg [(4'h8):(1'h0)] reg965 = (1'h0);
  reg [(3'h7):(1'h0)] reg964 = (1'h0);
  reg [(5'h14):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar962 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg961 = (1'h0);
  reg [(4'h9):(1'h0)] forvar960 = (1'h0);
  reg [(5'h12):(1'h0)] reg959 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg958 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg957 = (1'h0);
  reg [(3'h7):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar955 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg954 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg953 = (1'h0);
  reg signed [(4'he):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg951 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar950 = (1'h0);
  reg [(5'h12):(1'h0)] forvar949 = (1'h0);
  wire [(3'h6):(1'h0)] wire948;
  wire [(3'h7):(1'h0)] wire947;
  wire signed [(5'h14):(1'h0)] wire945;
  wire signed [(4'hf):(1'h0)] wire943;
  reg [(4'hc):(1'h0)] reg942 = (1'h0);
  reg [(5'h15):(1'h0)] reg941 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg938 = (1'h0);
  reg [(5'h13):(1'h0)] forvar937 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg936 = (1'h0);
  reg [(4'ha):(1'h0)] reg935 = (1'h0);
  reg [(4'ha):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar933 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg932 = (1'h0);
  wire [(2'h2):(1'h0)] wire931;
  wire [(4'hb):(1'h0)] wire929;
  wire [(4'he):(1'h0)] wire411;
  reg [(3'h5):(1'h0)] forvar5 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg7 = (1'h0);
  reg [(5'h10):(1'h0)] reg8 = (1'h0);
  reg [(5'h15):(1'h0)] reg9 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg10 = (1'h0);
  reg [(4'ha):(1'h0)] forvar11 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar12 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar14 = (1'h0);
  reg [(4'h8):(1'h0)] reg15 = (1'h0);
  reg [(3'h7):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg18 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg19 = (1'h0);
  reg [(5'h15):(1'h0)] reg20 = (1'h0);
  reg [(2'h2):(1'h0)] reg21 = (1'h0);
  reg [(3'h5):(1'h0)] forvar22 = (1'h0);
  reg [(2'h2):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar25 = (1'h0);
  reg [(4'h9):(1'h0)] reg26 = (1'h0);
  reg [(5'h14):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg28 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(5'h14):(1'h0)] forvar32 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg33 = (1'h0);
  reg signed [(4'he):(1'h0)] reg34 = (1'h0);
  reg [(4'h8):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar37 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar38 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg39 = (1'h0);
  reg [(4'hf):(1'h0)] forvar40 = (1'h0);
  reg [(3'h5):(1'h0)] reg41 = (1'h0);
  reg [(2'h3):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg43 = (1'h0);
  reg [(4'he):(1'h0)] reg44 = (1'h0);
  reg [(5'h10):(1'h0)] forvar45 = (1'h0);
  reg [(3'h7):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg47 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg49 = (1'h0);
  reg [(5'h15):(1'h0)] reg50 = (1'h0);
  reg [(5'h13):(1'h0)] reg51 = (1'h0);
  reg [(4'hd):(1'h0)] forvar52 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg53 = (1'h0);
  reg [(5'h12):(1'h0)] reg54 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg55 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg56 = (1'h0);
  reg [(4'hb):(1'h0)] reg57 = (1'h0);
  reg [(2'h3):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg59 = (1'h0);
  reg [(5'h15):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar61 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg62 = (1'h0);
  reg [(5'h15):(1'h0)] reg63 = (1'h0);
  reg [(5'h10):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg65 = (1'h0);
  reg [(4'hf):(1'h0)] reg66 = (1'h0);
  reg [(3'h5):(1'h0)] reg67 = (1'h0);
  reg [(3'h6):(1'h0)] reg68 = (1'h0);
  reg [(4'hc):(1'h0)] reg69 = (1'h0);
  reg [(5'h15):(1'h0)] reg70 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire409;
  assign y = {wire996,
                 reg995,
                 forvar994,
                 reg993,
                 reg986,
                 forvar984,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 forvar986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg979,
                 forvar978,
                 reg977,
                 forvar976,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 forvar969,
                 forvar968,
                 reg967,
                 forvar966,
                 reg965,
                 reg964,
                 reg963,
                 forvar962,
                 reg961,
                 forvar960,
                 reg959,
                 reg958,
                 reg957,
                 reg956,
                 forvar955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 forvar950,
                 forvar949,
                 wire948,
                 wire947,
                 wire945,
                 wire943,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg936,
                 reg935,
                 reg934,
                 forvar933,
                 reg932,
                 wire931,
                 wire929,
                 wire411,
                 forvar5,
                 forvar6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 forvar11,
                 forvar12,
                 reg13,
                 forvar14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 forvar22,
                 reg23,
                 reg24,
                 forvar25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 forvar32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 forvar37,
                 forvar38,
                 reg39,
                 forvar40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 forvar45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 forvar52,
                 reg53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 forvar60,
                 forvar61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 wire409,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar5 = (1'h0); (forvar5 < (2'h2)); forvar5 = (forvar5 + (1'h1)))
        begin
          for (forvar6 = (1'h0); (forvar6 < (2'h2)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 = (|(&$unsigned((wire2 | {forvar6}))));
              reg8 <= (forvar6[(1'h1):(1'h0)] ?
                  $signed(($unsigned(wire1[(3'h5):(3'h5)]) ?
                      $signed(reg7) : (~^wire3))) : wire3);
            end
          reg9 <= reg7[(4'h9):(3'h7)];
          reg10 <= ((8'ha3) || (~|$signed($unsigned((+forvar6)))));
        end
      for (forvar11 = (1'h0); (forvar11 < (2'h3)); forvar11 = (forvar11 + (1'h1)))
        begin
          for (forvar12 = (1'h0); (forvar12 < (2'h3)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 = (wire3[(1'h0):(1'h0)] ? $unsigned((8'h9d)) : (&wire0));
            end
          for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= $signed(forvar12[(3'h5):(3'h4)]);
              reg16 = reg8;
              reg17 = ($signed(wire0) ?
                  (wire1[(4'h8):(2'h2)] << $signed($signed($signed(reg15)))) : ($unsigned($signed(((8'hae) == reg8))) * {($signed(wire1) << $unsigned((8'hbf)))}));
              reg18 = wire4[(2'h3):(1'h0)];
              reg19 = (forvar11 ?
                  (+$unsigned(reg15[(2'h2):(2'h2)])) : (~&$signed((+$signed(reg13)))));
            end
        end
      reg20 = (7'h44);
      reg21 <= (wire2[(1'h1):(1'h0)] << (~&forvar12));
    end
  always
    @(posedge clk) begin
      for (forvar22 = (1'h0); (forvar22 < (2'h2)); forvar22 = (forvar22 + (1'h1)))
        begin
          if ((8'h9c))
            begin
              reg23 = $unsigned(($unsigned(reg7[(3'h5):(2'h2)]) * "XOLzsoZCLRT"));
            end
          else
            begin
              reg23 <= reg13[(4'hc):(4'h8)];
              reg24 <= wire2;
            end
          for (forvar25 = (1'h0); (forvar25 < (2'h3)); forvar25 = (forvar25 + (1'h1)))
            begin
              reg26 <= (($signed(reg21) != reg19) ? reg19 : forvar14);
              reg27 <= {(forvar25[(4'h9):(2'h3)] <<< $unsigned(("8h3JGe2mH" <= (forvar6 ?
                      reg13 : (8'ha2)))))};
              reg28 <= $signed(({($unsigned(wire3) ?
                      reg15[(4'h8):(3'h7)] : $unsigned(reg10))} <= ($signed((8'haf)) ?
                  reg10[(2'h3):(1'h1)] : (^(reg15 ? forvar6 : (8'hbf))))));
              reg29 <= reg8;
              reg30 <= $unsigned((((reg29 ? (-(8'ha3)) : {reg7, wire0}) ?
                      reg16[(3'h7):(1'h1)] : $signed($signed(forvar12))) ?
                  forvar12 : ($signed($signed(reg7)) > {$unsigned(reg27),
                      (reg27 >= (8'ha8))})));
            end
          reg31 <= (&forvar12);
          for (forvar32 = (1'h0); (forvar32 < (1'h1)); forvar32 = (forvar32 + (1'h1)))
            begin
              reg33 = (~|forvar25);
              reg34 = (forvar5[(1'h1):(1'h1)] ?
                  (~$signed((-(wire2 != forvar5)))) : ((^~$signed((^(8'ha6)))) & reg21[(1'h1):(1'h1)]));
            end
        end
      reg35 <= (($signed(wire2) + (8'hb6)) >>> {$unsigned(((reg30 >= reg33) ?
              ((8'hbc) ? reg24 : reg30) : (~|reg20)))});
      reg36 <= $unsigned($signed({$signed(reg13), reg15}));
      for (forvar37 = (1'h0); (forvar37 < (3'h4)); forvar37 = (forvar37 + (1'h1)))
        begin
          for (forvar38 = (1'h0); (forvar38 < (1'h0)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= $unsigned(reg17);
            end
          for (forvar40 = (1'h0); (forvar40 < (1'h0)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 <= $unsigned(((reg13 ?
                      (forvar37[(3'h4):(2'h3)] ?
                          (7'h44) : (reg36 ?
                              reg19 : reg23)) : "RRT1GsIryG94LHI") ?
                  forvar38 : $unsigned((reg15[(2'h2):(1'h1)] && (|reg34)))));
              reg42 <= {$unsigned((!{forvar14[(3'h6):(1'h0)], reg26})),
                  ((reg30 < (~^(forvar14 && (8'ha5)))) ?
                      ($unsigned((forvar37 ?
                          reg8 : reg19)) < reg35[(2'h3):(1'h1)]) : $unsigned(($signed(reg10) ?
                          $unsigned((8'ha7)) : (forvar22 & (8'ha8)))))};
            end
          reg43 <= ((^~reg7[(2'h2):(2'h2)]) >= ((($unsigned(reg41) ?
                      reg17[(4'ha):(1'h0)] : $unsigned(reg41)) ?
                  (|$signed(forvar40)) : $signed($unsigned(reg15))) ?
              (($unsigned(reg17) ? (reg18 ? (8'hae) : reg42) : forvar32) ?
                  forvar5 : (reg21[(1'h1):(1'h1)] | $signed(forvar12))) : {(wire3[(2'h2):(1'h1)] ?
                      $unsigned(reg33) : $signed(reg13)),
                  forvar38[(2'h2):(1'h0)]}));
          reg44 = wire2;
          for (forvar45 = (1'h0); (forvar45 < (1'h0)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 = (7'h40);
              reg47 = (~|($unsigned((8'hb2)) >> ((-(reg35 | forvar22)) ?
                  {(reg33 >= wire2)} : $signed(wire4[(4'ha):(2'h3)]))));
              reg48 <= forvar32[(3'h7):(1'h1)];
              reg49 <= forvar45;
              reg50 = (reg34 ?
                  (~|("" ?
                      $signed($signed(reg31)) : ((reg17 ~^ reg42) >> (~|forvar40)))) : "Qf9OCeSi9FZp9");
            end
        end
    end
  always
    @(posedge clk) begin
      reg51 <= ($signed($unsigned(reg7)) ?
          ((~^reg44[(4'h8):(1'h0)]) ~^ $unsigned((reg17[(4'h9):(3'h5)] ?
              $unsigned(reg47) : {reg27, forvar38}))) : forvar11);
      for (forvar52 = (1'h0); (forvar52 < (2'h2)); forvar52 = (forvar52 + (1'h1)))
        begin
          reg53 <= $signed(forvar5);
          if (($signed((|reg28[(5'h11):(4'hb)])) ?
              $unsigned($unsigned(((reg53 ? reg23 : (8'hbc)) ?
                  (reg53 > forvar5) : $signed((8'h9d))))) : reg8))
            begin
              reg54 <= reg43;
              reg55 = $unsigned((($signed((&forvar45)) ?
                  $signed((~^(8'ha3))) : $signed({forvar14})) ^ (((+(8'hbb)) != reg41) ?
                  ($unsigned(wire1) | $unsigned(forvar11)) : forvar37)));
              reg56 = (&$unsigned(reg24));
              reg57 <= (($unsigned((((7'h40) ? reg44 : (8'hb5)) ?
                      reg51[(4'h8):(3'h6)] : $signed(forvar11))) > ("" << {reg26,
                      (forvar32 > reg27)})) ?
                  ($unsigned($signed(reg26)) ?
                      $signed($unsigned({(7'h42)})) : (!reg35[(1'h1):(1'h0)])) : reg46[(1'h0):(1'h0)]);
            end
          else
            begin
              reg54 <= {$unsigned(forvar12), reg13};
              reg55 <= (forvar45[(3'h5):(2'h2)] ?
                  (!$signed((&(reg9 ? reg30 : (8'ha1))))) : reg57);
              reg56 <= (reg54[(2'h3):(1'h1)] ?
                  $signed($signed(($signed(reg8) ?
                      $signed(wire1) : (forvar5 - reg49)))) : reg57);
              reg57 <= ((^$signed(($signed((8'hbd)) ? (8'hba) : (^~reg26)))) ?
                  (reg20 & $signed(wire4)) : {((~|(reg41 ?
                              (8'h9f) : forvar11)) ?
                          $signed($unsigned(reg23)) : $signed((forvar5 - reg34)))});
              reg58 = (($signed({forvar14[(1'h1):(1'h0)], $signed(forvar6)}) ?
                  $unsigned((reg44 < forvar22[(3'h4):(2'h3)])) : reg29) >= ($signed((~^$unsigned(forvar45))) ?
                  ({(forvar52 ?
                          (8'hbc) : reg20)} == $unsigned($unsigned(reg57))) : reg31[(3'h7):(1'h1)]));
            end
        end
      reg59 <= $unsigned(reg54);
      for (forvar60 = (1'h0); (forvar60 < (2'h2)); forvar60 = (forvar60 + (1'h1)))
        begin
          for (forvar61 = (1'h0); (forvar61 < (1'h0)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 <= ({{wire0[(2'h2):(1'h0)]}} >= ({$signed(reg8),
                      ((forvar38 ? reg20 : forvar60) ^~ (~reg29))} ?
                  reg57 : (|(+(+reg23)))));
              reg63 <= reg23[(2'h2):(1'h0)];
              reg64 <= forvar22[(3'h4):(2'h3)];
              reg65 <= {({((~|reg31) ?
                          $signed(reg34) : $unsigned(forvar25))} & (reg18[(4'he):(4'h9)] || ((~&reg27) << reg57[(4'h8):(4'h8)]))),
                  $signed(wire2)};
              reg66 = (8'ha9);
            end
          if (reg16)
            begin
              reg67 <= ((($unsigned(((8'hbf) << reg20)) << $signed(reg58)) ?
                  ($signed($unsigned(forvar61)) ?
                      (~^$unsigned(reg28)) : wire3[(1'h1):(1'h0)]) : (($signed((8'hb9)) | reg57) ?
                      ($signed(reg20) ?
                          forvar61 : (wire4 ?
                              (8'had) : reg47)) : wire4)) == (!$signed(($unsigned(forvar14) - (reg23 >= reg66)))));
              reg68 <= ($unsigned($unsigned((forvar52 + (reg66 >> reg9)))) ?
                  reg20 : (-(~|($unsigned((8'hbc)) <= reg18))));
              reg69 <= reg36[(4'h9):(3'h5)];
              reg70 <= (reg66 < $signed({(((8'hb8) ?
                      reg46 : (8'hbb)) << (reg27 ? reg30 : forvar60)),
                  reg19}));
            end
          else
            begin
              reg67 <= (^~{$signed((reg66 > $unsigned(reg47)))});
              reg68 = {($signed({{forvar22}, (^(8'hbb))}) ?
                      $signed((8'hb3)) : forvar40[(4'ha):(3'h6)])};
              reg69 = $unsigned($signed(forvar40[(3'h4):(2'h3)]));
            end
        end
    end
  module71 modinst410 (wire409, clk, reg64, reg13, reg44, forvar52, reg66);
  assign wire411 = $signed((((-reg20[(3'h7):(2'h3)]) * forvar37) >= $signed(reg59[(1'h1):(1'h0)])));
  module412 modinst930 (.wire414(reg35), .wire416(reg68), .clk(clk), .wire413(reg8), .wire415(reg47), .y(wire929));
  assign wire931 = reg56;
  always
    @(posedge clk) begin
      reg932 <= (|((reg43 ?
          $signed($signed(reg59)) : (^wire2[(3'h7):(1'h1)])) << {$signed(forvar60),
          $unsigned((reg55 << reg18))}));
      for (forvar933 = (1'h0); (forvar933 < (2'h2)); forvar933 = (forvar933 + (1'h1)))
        begin
          if ((~&(|$unsigned((~|$unsigned(reg68))))))
            begin
              reg934 = $signed(((reg21 || (!{reg47, reg62})) ?
                  $unsigned(reg29) : (~|$unsigned(forvar6[(2'h2):(2'h2)]))));
              reg935 = $unsigned($unsigned((($signed(forvar61) << $signed(reg35)) ?
                  (^~(reg24 ? wire2 : reg36)) : reg10)));
              reg936 = reg34[(2'h2):(2'h2)];
            end
          else
            begin
              reg934 = (~&(^~"aSltyDBf"));
              reg935 = (($signed(reg17[(4'h9):(3'h6)]) ?
                      ($unsigned(forvar6) ?
                          $unsigned($unsigned(reg34)) : $unsigned((wire411 ?
                              (8'haf) : reg24))) : (reg54 ?
                          forvar14 : (wire1 ?
                              (reg39 ?
                                  (8'h9f) : reg35) : forvar5[(2'h2):(2'h2)]))) ?
                  wire0[(4'hf):(4'h9)] : {$signed($unsigned((forvar61 == forvar12))),
                      wire929[(4'hb):(3'h5)]});
            end
          for (forvar937 = (1'h0); (forvar937 < (1'h0)); forvar937 = (forvar937 + (1'h1)))
            begin
              reg938 <= (-("bdnRUXkRJVbvAs2R" ?
                  (~|($unsigned((8'hb7)) == $signed(reg50))) : "TTUl"));
              reg939 <= (^~wire4);
              reg940 = reg17[(2'h2):(1'h1)];
              reg941 <= $unsigned(reg24);
              reg942 = ((($unsigned($unsigned(reg936)) ?
                      (!(reg66 >> reg51)) : ($signed((8'hb8)) ?
                          ((8'ha5) ^~ reg939) : (wire4 == reg19))) ?
                  ({(^reg932)} ?
                      reg24[(4'hd):(2'h3)] : (&{(8'hb0),
                          reg15})) : {"VqUtqrUzSWg6oaWxuDKb",
                      $unsigned("5VqEh2WDw2Sy")}) ^ ($signed(reg30[(4'hf):(4'ha)]) ?
                  (forvar52 > ("" | $unsigned((8'ha8)))) : ($signed(forvar937[(4'hd):(4'h9)]) <<< wire2)));
            end
        end
    end
  module832 modinst944 (.clk(clk), .y(wire943), .wire836(reg9), .wire834(reg51), .wire835(reg36), .wire833(reg935));
  module442 modinst946 (.y(wire945), .wire444(reg70), .wire443(reg934), .wire445(wire4), .wire446(reg938), .clk(clk));
  assign wire947 = ($signed($signed($signed((wire0 || (8'ha8))))) || reg23);
  assign wire948 = $signed($signed(((!$unsigned(reg13)) | ({(8'hba), forvar37} ?
                       $unsigned(reg938) : {forvar5, reg64}))));
  always
    @(posedge clk) begin
      for (forvar949 = (1'h0); (forvar949 < (2'h2)); forvar949 = (forvar949 + (1'h1)))
        begin
          for (forvar950 = (1'h0); (forvar950 < (3'h4)); forvar950 = (forvar950 + (1'h1)))
            begin
              reg951 = reg44[(2'h3):(2'h2)];
              reg952 = reg51[(2'h2):(2'h2)];
              reg953 <= forvar45;
              reg954 = $unsigned("bsmJrNyEUSulgo9dQsXB");
            end
          for (forvar955 = (1'h0); (forvar955 < (1'h0)); forvar955 = (forvar955 + (1'h1)))
            begin
              reg956 = wire3[(2'h3):(1'h0)];
              reg957 <= reg956[(1'h0):(1'h0)];
              reg958 <= (&($signed((reg942[(2'h2):(1'h1)] << (reg64 != (7'h44)))) ?
                  $unsigned({$unsigned(wire947),
                      $unsigned(reg29)}) : (({forvar40} && $signed(reg57)) ?
                      ({reg70} + $unsigned(reg43)) : forvar6)));
              reg959 = reg952[(2'h2):(2'h2)];
            end
          for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
            begin
              reg961 = {(^~$signed(((reg34 == forvar60) ?
                      (reg68 & reg26) : $signed(wire2)))),
                  (+$signed(forvar937[(4'hc):(3'h5)]))};
            end
          for (forvar962 = (1'h0); (forvar962 < (2'h3)); forvar962 = (forvar962 + (1'h1)))
            begin
              reg963 <= $signed({forvar12[(1'h0):(1'h0)],
                  "KHGz2gMeXBJntqpc2i"});
              reg964 = reg28[(3'h7):(3'h5)];
              reg965 = reg58[(1'h1):(1'h0)];
            end
          for (forvar966 = (1'h0); (forvar966 < (2'h3)); forvar966 = (forvar966 + (1'h1)))
            begin
              reg967 <= ((~&($signed((reg959 != reg70)) ?
                      ((wire929 ?
                          forvar937 : reg935) ~^ $unsigned(reg8)) : $unsigned({reg70,
                          (8'hb2)}))) ?
                  {((reg16 ? (8'h9e) : reg18[(3'h6):(1'h1)]) ?
                          ((reg31 ^ reg51) ?
                              (reg942 ?
                                  wire3 : (8'hbb)) : (+forvar950)) : ($signed((7'h43)) << {forvar40})),
                      ($signed((wire0 ? (8'ha8) : reg961)) ?
                          (~|$signed(reg9)) : "ol")} : $signed(reg33[(2'h2):(1'h1)]));
            end
        end
      for (forvar968 = (1'h0); (forvar968 < (1'h1)); forvar968 = (forvar968 + (1'h1)))
        begin
          for (forvar969 = (1'h0); (forvar969 < (1'h1)); forvar969 = (forvar969 + (1'h1)))
            begin
              reg970 <= ({$unsigned(reg935[(3'h7):(3'h4)])} ?
                  {$unsigned(forvar52)} : reg48);
              reg971 <= ($unsigned(("1ssooU0uQ" ^~ (8'hb1))) ?
                  $unsigned((~^{{forvar52}})) : (forvar22[(2'h2):(2'h2)] <= reg65[(2'h2):(2'h2)]));
              reg972 <= ($signed({(8'hba)}) ?
                  $unsigned($unsigned($unsigned(wire948[(3'h4):(1'h1)]))) : ({$signed((reg957 ^ wire945)),
                          $signed("IZXUOIlex9pBZqdpEO")} ?
                      $signed(({reg941,
                          reg20} << $signed(wire929))) : wire947[(3'h4):(1'h0)]));
              reg973 <= $signed(wire929);
              reg974 <= ((((reg65 * $signed(reg28)) & $signed({reg942,
                      (7'h40)})) ?
                  ((8'hbd) & $unsigned((reg48 ?
                      reg29 : forvar45))) : $unsigned((wire945 | (forvar968 && reg41)))) * reg10);
            end
          reg975 <= reg26[(4'h8):(3'h6)];
          for (forvar976 = (1'h0); (forvar976 < (2'h3)); forvar976 = (forvar976 + (1'h1)))
            begin
              reg977 = (~&$unsigned("v7BDkN"));
            end
          for (forvar978 = (1'h0); (forvar978 < (1'h1)); forvar978 = (forvar978 + (1'h1)))
            begin
              reg979 <= $unsigned((({$signed((8'h9f)),
                      (reg69 << reg951)} && reg64) ?
                  {reg16,
                      $signed($signed(reg44))} : (($signed(reg952) && (7'h41)) <<< $unsigned(reg68[(1'h0):(1'h0)]))));
              reg980 = wire943[(4'hb):(4'ha)];
              reg981 <= $unsigned($signed({(-$unsigned(forvar949))}));
              reg982 = forvar933[(1'h1):(1'h0)];
            end
          reg983 <= (wire409 ?
              (~$unsigned("viDtXRVtUnkqCb")) : $unsigned(((reg958 ?
                  "9amz2" : $unsigned(reg34)) >>> "gH")));
        end
      if ($unsigned($signed($unsigned(((+wire945) ?
          (forvar22 ? wire3 : (8'hb7)) : forvar950)))))
        begin
          if (reg67)
            begin
              reg984 <= $signed(((-reg50[(1'h1):(1'h0)]) ?
                  $signed((forvar38 || $unsigned(reg39))) : reg942));
              reg985 <= (~^wire4[(4'h9):(3'h7)]);
            end
          else
            begin
              reg984 <= (wire948 << $unsigned((reg33 <<< (8'ha0))));
            end
          for (forvar986 = (1'h0); (forvar986 < (1'h0)); forvar986 = (forvar986 + (1'h1)))
            begin
              reg987 <= ((reg938 == reg941[(4'h9):(2'h3)]) ?
                  $signed("RksiF6oiRJ0Y") : (|{$unsigned(reg21[(2'h2):(1'h1)])}));
              reg988 <= forvar37[(2'h3):(1'h1)];
              reg989 <= forvar986[(3'h5):(2'h3)];
            end
          if (reg66[(3'h5):(1'h0)])
            begin
              reg990 <= (&$signed((reg30 ?
                  forvar968 : {(reg940 ? wire409 : forvar966), (!wire947)})));
              reg991 = $signed($unsigned((^($unsigned((8'hbc)) > {wire4}))));
            end
          else
            begin
              reg990 = $signed($unsigned($unsigned(("" >> (-reg23)))));
              reg991 = $unsigned($unsigned($unsigned((forvar6 ?
                  reg964[(2'h3):(1'h1)] : (reg956 <<< reg63)))));
              reg992 <= {(~(^~$signed(((8'hb3) ? reg68 : reg965)))),
                  $signed($signed(forvar986))};
            end
        end
      else
        begin
          for (forvar984 = (1'h0); (forvar984 < (2'h3)); forvar984 = (forvar984 + (1'h1)))
            begin
              reg985 = $signed("h03NXa3kbhplgsW8Tc2p");
              reg986 <= (wire945 ?
                  $signed($signed(((~(8'hbc)) ?
                      (~wire411) : (~reg57)))) : (wire948[(3'h4):(1'h1)] >= (!$signed((reg54 ?
                      reg939 : reg970)))));
              reg987 = "4XIVgltP8WI7gm6CK";
            end
          if (wire3)
            begin
              reg988 <= $unsigned($signed(forvar986));
              reg989 = (~$signed($signed($signed((^reg932)))));
              reg990 = reg989;
            end
          else
            begin
              reg988 <= reg9;
              reg989 = forvar25[(5'h12):(3'h5)];
              reg990 <= "W5oWd3nxQs2TVZiU";
              reg991 <= (-(&reg984[(4'h9):(4'h8)]));
            end
        end
      reg993 = reg15;
      for (forvar994 = (1'h0); (forvar994 < (1'h1)); forvar994 = (forvar994 + (1'h1)))
        begin
          reg995 <= (8'hb7);
        end
    end
  assign wire996 = reg967[(3'h7):(3'h7)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module412  (y, clk, wire416, wire415, wire414, wire413);
  output wire [(32'h5f7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire416;
  input wire signed [(3'h7):(1'h0)] wire415;
  input wire [(4'h8):(1'h0)] wire414;
  input wire signed [(3'h5):(1'h0)] wire413;
  wire signed [(2'h2):(1'h0)] wire928;
  wire signed [(5'h13):(1'h0)] wire926;
  wire signed [(5'h12):(1'h0)] wire831;
  wire [(4'h9):(1'h0)] wire830;
  wire [(4'h9):(1'h0)] wire829;
  wire [(4'h9):(1'h0)] wire828;
  reg signed [(4'ha):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg826 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg825 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg824 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg823 = (1'h0);
  reg [(4'hd):(1'h0)] reg822 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg821 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar820 = (1'h0);
  reg [(4'hc):(1'h0)] forvar819 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg818 = (1'h0);
  reg [(4'h9):(1'h0)] reg817 = (1'h0);
  reg [(5'h13):(1'h0)] reg816 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg815 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg814 = (1'h0);
  reg [(3'h4):(1'h0)] reg813 = (1'h0);
  reg [(3'h6):(1'h0)] forvar812 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg811 = (1'h0);
  reg [(3'h6):(1'h0)] reg810 = (1'h0);
  reg signed [(4'he):(1'h0)] reg809 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg808 = (1'h0);
  reg [(5'h12):(1'h0)] reg807 = (1'h0);
  reg [(5'h11):(1'h0)] forvar806 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire805;
  reg signed [(3'h5):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg802 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg801 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg800 = (1'h0);
  reg [(4'hf):(1'h0)] forvar799 = (1'h0);
  reg [(5'h10):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg797 = (1'h0);
  reg [(3'h4):(1'h0)] reg796 = (1'h0);
  reg [(5'h11):(1'h0)] forvar795 = (1'h0);
  reg [(4'hc):(1'h0)] forvar794 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg781 = (1'h0);
  reg [(3'h5):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg792 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg791 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg790 = (1'h0);
  reg [(5'h10):(1'h0)] forvar789 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg788 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg787 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg786 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg785 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg784 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg783 = (1'h0);
  reg [(3'h6):(1'h0)] reg782 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar781 = (1'h0);
  reg [(3'h6):(1'h0)] reg780 = (1'h0);
  reg [(4'hb):(1'h0)] reg779 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar778 = (1'h0);
  reg [(4'ha):(1'h0)] reg777 = (1'h0);
  reg [(5'h10):(1'h0)] reg776 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire775;
  reg signed [(2'h3):(1'h0)] reg774 = (1'h0);
  reg [(4'h8):(1'h0)] reg773 = (1'h0);
  reg [(5'h13):(1'h0)] reg772 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar771 = (1'h0);
  reg [(4'ha):(1'h0)] reg770 = (1'h0);
  reg [(5'h11):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg768 = (1'h0);
  reg [(4'hb):(1'h0)] reg767 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar766 = (1'h0);
  reg [(4'hb):(1'h0)] reg765 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg764 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg763 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg762 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg761 = (1'h0);
  reg [(3'h7):(1'h0)] reg760 = (1'h0);
  reg [(3'h6):(1'h0)] forvar759 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar758 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg757 = (1'h0);
  reg [(4'hb):(1'h0)] reg756 = (1'h0);
  reg [(3'h6):(1'h0)] reg755 = (1'h0);
  reg [(4'hd):(1'h0)] reg754 = (1'h0);
  reg [(5'h14):(1'h0)] forvar753 = (1'h0);
  reg [(5'h14):(1'h0)] reg752 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg751 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg750 = (1'h0);
  reg [(2'h2):(1'h0)] reg749 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg747 = (1'h0);
  reg [(4'he):(1'h0)] reg746 = (1'h0);
  reg [(4'he):(1'h0)] reg745 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar744 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg743 = (1'h0);
  reg [(4'hf):(1'h0)] reg742 = (1'h0);
  reg [(5'h11):(1'h0)] forvar741 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg740 = (1'h0);
  reg [(4'he):(1'h0)] reg739 = (1'h0);
  reg [(5'h13):(1'h0)] reg738 = (1'h0);
  reg [(4'he):(1'h0)] reg737 = (1'h0);
  reg [(4'h9):(1'h0)] reg736 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar735 = (1'h0);
  reg [(4'h8):(1'h0)] forvar734 = (1'h0);
  reg [(4'hd):(1'h0)] reg733 = (1'h0);
  wire [(4'h8):(1'h0)] wire731;
  wire [(5'h14):(1'h0)] wire643;
  wire [(5'h13):(1'h0)] wire441;
  reg signed [(2'h3):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg439 = (1'h0);
  reg [(5'h12):(1'h0)] forvar438 = (1'h0);
  reg [(4'ha):(1'h0)] reg437 = (1'h0);
  reg [(4'hb):(1'h0)] reg436 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar435 = (1'h0);
  wire [(4'ha):(1'h0)] wire434;
  reg signed [(5'h15):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg432 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg431 = (1'h0);
  reg [(4'h9):(1'h0)] reg430 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg429 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar427 = (1'h0);
  reg [(3'h7):(1'h0)] reg426 = (1'h0);
  reg [(5'h11):(1'h0)] reg425 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg424 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar423 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar422 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg421 = (1'h0);
  reg [(5'h15):(1'h0)] reg420 = (1'h0);
  reg [(5'h10):(1'h0)] reg419 = (1'h0);
  wire [(4'ha):(1'h0)] wire418;
  wire [(5'h13):(1'h0)] wire417;
  assign y = {wire928,
                 wire926,
                 wire831,
                 wire830,
                 wire829,
                 wire828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 forvar820,
                 forvar819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 forvar812,
                 reg811,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 forvar806,
                 wire805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 forvar799,
                 reg798,
                 reg797,
                 reg796,
                 forvar795,
                 forvar794,
                 reg781,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 forvar789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 forvar781,
                 reg780,
                 reg779,
                 forvar778,
                 reg777,
                 reg776,
                 wire775,
                 reg774,
                 reg773,
                 reg772,
                 forvar771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 forvar766,
                 reg765,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg760,
                 forvar759,
                 forvar758,
                 reg757,
                 reg756,
                 reg755,
                 reg754,
                 forvar753,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 forvar744,
                 reg743,
                 reg742,
                 forvar741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 forvar735,
                 forvar734,
                 reg733,
                 wire731,
                 wire643,
                 wire441,
                 reg440,
                 reg439,
                 forvar438,
                 reg437,
                 reg436,
                 forvar435,
                 wire434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 reg426,
                 reg425,
                 reg424,
                 forvar423,
                 forvar422,
                 reg421,
                 reg420,
                 reg419,
                 wire418,
                 wire417,
                 (1'h0)};
  assign wire417 = wire415;
  assign wire418 = wire417[(4'hf):(4'hc)];
  always
    @(posedge clk) begin
      reg419 <= (wire415[(1'h1):(1'h0)] ?
          {wire413[(2'h3):(2'h2)]} : ($unsigned("kPLOR751") >> {$unsigned($signed(wire417)),
              $unsigned((~^wire414))}));
      reg420 = ((($unsigned(wire414) ?
              $unsigned(wire416[(2'h3):(1'h1)]) : (wire416[(3'h4):(3'h4)] ^~ (wire415 != reg419))) ?
          wire415 : wire417) - (~^(wire413 ?
          wire414[(3'h6):(2'h2)] : $unsigned({reg419, wire415}))));
      reg421 <= (|{(-$signed({wire418}))});
      for (forvar422 = (1'h0); (forvar422 < (2'h3)); forvar422 = (forvar422 + (1'h1)))
        begin
          for (forvar423 = (1'h0); (forvar423 < (2'h2)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 <= reg420;
              reg425 <= (~&$signed((((&reg419) ?
                  wire417 : $unsigned(wire418)) >>> $signed(reg420[(2'h3):(2'h3)]))));
              reg426 <= (($unsigned(((+forvar423) ?
                  $unsigned(reg419) : {(8'ha3),
                      wire417})) & forvar422) > ($signed($unsigned($signed(reg419))) ?
                  ("9gfdN7akAOA1Zxks" ?
                      "p7LLEC18" : wire418[(4'h8):(3'h6)]) : ({{(8'ha2),
                          (8'hb3)}} == $signed(wire413[(1'h1):(1'h1)]))));
            end
          for (forvar427 = (1'h0); (forvar427 < (2'h3)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= ($signed(((~|$signed((7'h42))) * wire413[(2'h3):(2'h3)])) ?
                  $unsigned((|wire415)) : ((-wire413) ?
                      ($unsigned(reg424) << $signed((reg425 >> wire417))) : $signed(((wire413 ?
                              (8'hb7) : forvar423) ?
                          (wire416 >>> wire414) : (reg420 ?
                              reg421 : reg424)))));
              reg429 <= (reg425[(4'ha):(2'h3)] ?
                  (~|wire416[(3'h4):(1'h1)]) : $signed($unsigned(({reg428} ?
                      reg425 : (^(8'hba))))));
              reg430 <= (({({reg429, wire415} ?
                              forvar422[(4'hd):(4'hc)] : reg425),
                          $unsigned($unsigned(wire417))} ?
                      (+forvar422[(3'h7):(3'h4)]) : wire414[(1'h0):(1'h0)]) ?
                  (reg429 ?
                      wire417[(1'h1):(1'h0)] : ({$signed(reg425),
                          wire415[(2'h3):(2'h3)]} ^ (~&(reg424 == wire416)))) : ({reg419} < (reg419[(4'he):(2'h2)] ?
                      $unsigned(wire413) : ($unsigned(wire413) ?
                          reg420 : $unsigned(reg419)))));
              reg431 <= ((wire413 ?
                      wire413[(1'h0):(1'h0)] : {$signed((forvar427 ?
                              reg419 : wire415))}) ?
                  ((reg430 ?
                      $signed($signed((8'hbc))) : ($signed(wire416) >> $unsigned(forvar423))) || $unsigned(wire414)) : (+(8'hb3)));
            end
          reg432 <= reg426;
        end
      reg433 = {"RvOHg",
          (($signed($signed(reg426)) ?
              {((8'hb2) << (7'h42)),
                  reg432[(1'h0):(1'h0)]} : ($signed((8'hac)) ?
                  {wire416, reg429} : (-wire417))) == ({(!wire413)} ?
              $unsigned((reg432 ? reg432 : wire417)) : (!$signed(wire418))))};
    end
  assign wire434 = reg420;
  always
    @(posedge clk) begin
      for (forvar435 = (1'h0); (forvar435 < (2'h2)); forvar435 = (forvar435 + (1'h1)))
        begin
          reg436 = (!($signed(forvar423) * $signed({{reg430, wire413},
              (reg429 >> reg425)})));
          reg437 = (-reg429);
          for (forvar438 = (1'h0); (forvar438 < (1'h1)); forvar438 = (forvar438 + (1'h1)))
            begin
              reg439 = (((((wire415 ? reg436 : reg429) ?
                      (forvar423 && reg428) : "9QCW69UezUR") - {((8'hbb) ?
                          (7'h44) : forvar435)}) ?
                  (8'ha0) : ((&(wire413 & (8'hb1))) <= reg430[(1'h1):(1'h1)])) + ($signed((((7'h41) ?
                          (8'hbd) : reg426) ?
                      (8'ha5) : wire434)) ?
                  (($signed(wire413) ?
                      $unsigned(wire417) : (wire415 ?
                          forvar422 : (8'hb5))) - (~|(reg433 + reg431))) : (~&$unsigned($unsigned(wire434)))));
              reg440 <= {(reg432[(4'hc):(2'h2)] ?
                      ($unsigned(wire413) ?
                          wire417[(4'ha):(2'h3)] : $unsigned(reg439)) : (wire418[(3'h4):(3'h4)] ?
                          reg421 : (|((8'hbf) ? reg431 : wire413)))),
                  $signed({(+$signed((8'hb1)))})};
            end
        end
    end
  assign wire441 = (~forvar423);
  module442 modinst644 (.clk(clk), .y(wire643), .wire444(reg420), .wire445(wire415), .wire446(wire413), .wire443(reg425));
  module645 modinst732 (.wire649(wire441), .y(wire731), .clk(clk), .wire647(reg430), .wire648(forvar427), .wire646(reg432));
  always
    @(posedge clk) begin
      reg733 <= $unsigned((reg425 ?
          ($signed((^~reg424)) ^ forvar423) : $unsigned("kB")));
      for (forvar734 = (1'h0); (forvar734 < (2'h2)); forvar734 = (forvar734 + (1'h1)))
        begin
          for (forvar735 = (1'h0); (forvar735 < (1'h0)); forvar735 = (forvar735 + (1'h1)))
            begin
              reg736 <= (wire414[(1'h0):(1'h0)] >= reg430[(1'h0):(1'h0)]);
              reg737 <= wire418[(3'h7):(1'h0)];
              reg738 <= reg429;
              reg739 <= ($signed(($unsigned((|wire416)) == $unsigned(reg428))) < $signed(({$unsigned(reg419),
                      reg431[(3'h5):(1'h1)]} ?
                  $unsigned((~&forvar423)) : reg738)));
            end
          reg740 = reg738[(4'h8):(1'h0)];
          for (forvar741 = (1'h0); (forvar741 < (1'h0)); forvar741 = (forvar741 + (1'h1)))
            begin
              reg742 <= {{$signed(forvar734[(2'h2):(1'h1)])},
                  ($signed({$signed(wire417)}) ?
                      $unsigned(reg439) : (reg738[(2'h3):(1'h1)] ?
                          $signed(reg421[(4'hc):(1'h0)]) : $unsigned({reg739})))};
            end
        end
      reg743 <= forvar435;
      if (forvar734[(2'h2):(1'h1)])
        begin
          for (forvar744 = (1'h0); (forvar744 < (1'h0)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= ("bK1Yx1DFxsd" >>> (forvar735[(1'h1):(1'h0)] ?
                  (+reg420) : {$unsigned($unsigned((8'ha6))),
                      ($unsigned(forvar427) ^~ (reg740 ? (7'h43) : wire416))}));
              reg746 = (reg433 ~^ ({reg433, {{reg437, wire441}}} ?
                  $unsigned((~|$unsigned(forvar741))) : $unsigned(reg425)));
              reg747 <= wire413[(3'h5):(3'h4)];
            end
        end
      else
        begin
          for (forvar744 = (1'h0); (forvar744 < (1'h0)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= $signed(($signed({(reg739 >= reg440), reg436}) ?
                  (7'h42) : reg429[(4'hd):(4'ha)]));
              reg746 = (-forvar741);
              reg747 <= (((reg429 << {$signed(forvar734),
                      reg739[(2'h2):(2'h2)]}) && $unsigned((8'hbd))) ?
                  (~|($unsigned($unsigned(reg421)) ?
                      {reg440, wire416} : ((wire416 ?
                          reg440 : reg439) & ((8'ha4) ?
                          reg740 : reg421)))) : {"wNw"});
              reg748 = reg426;
              reg749 = wire414;
            end
          reg750 <= {reg437[(3'h4):(3'h4)]};
        end
      reg751 <= ((($signed((^~reg742)) >> $signed($unsigned(reg740))) ?
              {$signed($unsigned((7'h40))),
                  ($unsigned(wire441) ?
                      (-reg424) : reg745[(4'h9):(3'h5)])} : reg733[(4'h9):(2'h2)]) ?
          $signed(reg745) : {{$signed(wire414[(3'h4):(1'h0)])}});
    end
  always
    @(posedge clk) begin
      reg752 <= reg429[(4'ha):(4'h9)];
      for (forvar753 = (1'h0); (forvar753 < (3'h4)); forvar753 = (forvar753 + (1'h1)))
        begin
          reg754 <= (reg440[(1'h0):(1'h0)] ?
              $signed(forvar735[(3'h4):(3'h4)]) : reg420);
          reg755 <= wire413[(1'h0):(1'h0)];
          reg756 <= reg437;
          reg757 = (&((((7'h41) * (wire731 ? reg742 : wire415)) ?
              ((reg440 <= reg740) >>> reg425) : $unsigned((reg425 && reg436))) ^~ reg428[(1'h1):(1'h0)]));
        end
      for (forvar758 = (1'h0); (forvar758 < (2'h3)); forvar758 = (forvar758 + (1'h1)))
        begin
          for (forvar759 = (1'h0); (forvar759 < (1'h0)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 <= $signed(((~^(wire731[(3'h4):(1'h0)] & (+reg431))) ?
                  reg439 : (^$unsigned($unsigned(wire417)))));
              reg761 <= $unsigned($unsigned(reg751[(2'h3):(1'h0)]));
            end
          reg762 <= ($signed(((reg430 ?
                  $signed((8'ha8)) : (reg733 ? wire417 : wire643)) ?
              reg756[(3'h7):(2'h2)] : (&reg740[(3'h5):(1'h0)]))) >>> ("gyKFtbXPte" > {$signed(reg433[(3'h7):(1'h1)]),
              ((reg433 ? reg754 : forvar422) ?
                  {reg756} : reg761[(2'h2):(1'h1)])}));
          if ($unsigned({(reg736[(3'h4):(2'h2)] ?
                  wire417 : {$unsigned(reg756), (reg748 * forvar744)})}))
            begin
              reg763 <= reg425;
              reg764 <= {{reg737[(4'hb):(4'ha)],
                      $signed(((~^(7'h41)) <= (reg431 - reg762)))}};
              reg765 = reg430;
            end
          else
            begin
              reg763 <= reg738;
            end
          for (forvar766 = (1'h0); (forvar766 < (2'h2)); forvar766 = (forvar766 + (1'h1)))
            begin
              reg767 = ($signed({reg748}) || (reg756[(3'h7):(3'h4)] ?
                  (((!reg440) ?
                      (forvar741 ?
                          (8'hb8) : forvar435) : reg739[(4'hb):(3'h5)]) && (wire434 && (8'hb3))) : reg426[(3'h7):(3'h5)]));
              reg768 <= (~&(8'h9d));
              reg769 <= (^($signed(((^forvar435) >= $unsigned(reg425))) && reg749));
              reg770 = forvar758[(3'h7):(2'h3)];
            end
          for (forvar771 = (1'h0); (forvar771 < (2'h3)); forvar771 = (forvar771 + (1'h1)))
            begin
              reg772 <= (wire434[(3'h7):(3'h7)] ?
                  $signed((8'hb7)) : $unsigned(reg755));
              reg773 = (~^wire643);
            end
        end
      reg774 = $signed((~$unsigned(((reg762 > reg761) == (+(8'hb2))))));
    end
  assign wire775 = wire441[(3'h6):(2'h3)];
  always
    @(posedge clk) begin
      reg776 = ({$signed((((8'ha9) ? reg428 : reg751) + reg761[(2'h3):(1'h0)])),
          reg755[(2'h2):(2'h2)]} ^~ $unsigned($unsigned("G0FrpncHpLGhmd0y")));
      reg777 = (^forvar741);
      for (forvar778 = (1'h0); (forvar778 < (2'h2)); forvar778 = (forvar778 + (1'h1)))
        begin
          reg779 <= reg426;
          reg780 <= $unsigned(((~reg754) << (-$signed(reg743[(5'h10):(4'hf)]))));
        end
      if ($unsigned((^(8'hac))))
        begin
          for (forvar781 = (1'h0); (forvar781 < (2'h3)); forvar781 = (forvar781 + (1'h1)))
            begin
              reg782 <= (({(^{reg431, wire415}),
                      $unsigned((|reg420))} != ((forvar759 ?
                          {reg421} : (&reg761)) ?
                      $unsigned("hcUULVLeGFY") : forvar753)) ?
                  forvar734 : (~|wire731));
            end
          reg783 <= $signed(wire731[(3'h6):(2'h2)]);
          if (((((^(reg737 <<< reg765)) ?
              {$unsigned((8'hb2)),
                  reg425} : $unsigned(reg742)) >> reg740) < (8'hba)))
            begin
              reg784 <= (reg430[(3'h5):(2'h3)] ?
                  $unsigned($signed($signed($unsigned(reg424)))) : reg770);
            end
          else
            begin
              reg784 <= (-forvar744);
              reg785 = ($signed(((reg747 ? $signed(reg742) : (^reg433)) ?
                  reg749[(1'h1):(1'h0)] : {$signed(reg437)})) > wire731);
              reg786 <= (8'hb6);
              reg787 <= (~&("JtgkAVtvS" + ((reg436 ?
                  reg426[(3'h5):(2'h2)] : (reg764 ?
                      forvar744 : wire414)) | (8'ha6))));
              reg788 <= "24FGAxtrpA";
            end
          for (forvar789 = (1'h0); (forvar789 < (3'h4)); forvar789 = (forvar789 + (1'h1)))
            begin
              reg790 <= {(8'h9f), reg762};
              reg791 <= (|($signed((7'h42)) | ((~^(forvar771 - (8'hb0))) & $signed({forvar735,
                  reg790}))));
              reg792 <= ("38wF1zftRJMUb" | (reg745 < (($unsigned((8'hb7)) + $signed(reg772)) < (wire434 << (~|(8'ha7))))));
              reg793 = ((|forvar758[(3'h7):(1'h0)]) & forvar734);
            end
        end
      else
        begin
          if ($unsigned($signed($signed((~&(~reg755))))))
            begin
              reg781 <= reg742;
              reg782 <= reg784[(3'h7):(2'h3)];
              reg783 = $unsigned(reg747);
            end
          else
            begin
              reg781 = (forvar766[(4'hd):(3'h4)] >>> ("TB2d" << $signed(($signed(forvar778) != ((8'had) <= reg786)))));
            end
          if (($unsigned((((reg432 ^ reg420) ^ reg745) <= reg430)) + ((((reg755 < reg733) ?
              {reg761} : (8'ha1)) ~^ $signed((reg428 ?
              forvar435 : wire441))) * (((8'hb4) ?
                  $unsigned(reg739) : (8'hb7)) ?
              reg793 : ({(8'hab), (8'ha1)} ? (reg792 + reg783) : (!reg431))))))
            begin
              reg784 <= ($signed((forvar741[(4'h8):(2'h2)] ?
                      ($signed(reg429) <<< reg740) : (+$signed(reg431)))) ?
                  {$signed((reg432 >> (reg792 ?
                          reg430 : reg752)))} : (~|$signed($signed(wire643))));
              reg785 <= $signed($signed((~|$signed($signed(forvar744)))));
              reg786 <= ($unsigned((~^reg777[(3'h4):(1'h0)])) >>> (reg779[(4'hb):(3'h7)] ?
                  reg437 : (^~($unsigned(wire416) ?
                      forvar789 : $signed(reg774)))));
              reg787 <= $signed($signed((reg770[(3'h6):(1'h0)] ?
                  forvar781 : (|(reg751 ? reg767 : reg433)))));
              reg788 <= $unsigned(reg425[(4'h8):(3'h6)]);
            end
          else
            begin
              reg784 = reg762;
              reg785 = (forvar427 - (|reg421[(5'h11):(3'h4)]));
              reg786 <= reg432[(3'h7):(3'h4)];
              reg787 <= {(!($unsigned(reg793) ?
                      $unsigned((reg791 ?
                          reg768 : reg742)) : $signed((reg439 != reg437))))};
              reg788 <= (8'hbe);
            end
        end
      for (forvar794 = (1'h0); (forvar794 < (1'h0)); forvar794 = (forvar794 + (1'h1)))
        begin
          for (forvar795 = (1'h0); (forvar795 < (2'h3)); forvar795 = (forvar795 + (1'h1)))
            begin
              reg796 = (((&reg783) ?
                  $signed(reg783[(2'h2):(2'h2)]) : $unsigned((reg436 ?
                      (~reg760) : $unsigned(reg742)))) ~^ ($unsigned((8'h9e)) ?
                  {reg740[(2'h2):(1'h1)], reg751} : (~&(((8'ha3) ?
                      reg792 : (7'h42)) - (reg764 ? reg754 : reg764)))));
              reg797 <= $unsigned(reg421);
              reg798 <= ({$signed((~^(wire775 == forvar789))),
                  (reg756 | (~|$unsigned(wire414)))} >> ((!reg784[(2'h2):(1'h1)]) & $unsigned(reg756)));
            end
          for (forvar799 = (1'h0); (forvar799 < (2'h3)); forvar799 = (forvar799 + (1'h1)))
            begin
              reg800 = (wire418 >= $signed($signed(((+forvar758) ~^ $signed(reg755)))));
              reg801 = ({{(forvar427 ?
                              (reg767 ? reg787 : wire413) : (wire418 ?
                                  reg798 : reg791))}} ?
                  reg756[(2'h3):(2'h3)] : $unsigned((&$unsigned((reg439 * wire416)))));
            end
          reg802 <= reg740;
          reg803 = reg762[(3'h5):(3'h5)];
          reg804 <= reg772[(5'h13):(1'h0)];
        end
    end
  assign wire805 = reg785;
  always
    @(posedge clk) begin
      for (forvar806 = (1'h0); (forvar806 < (1'h1)); forvar806 = (forvar806 + (1'h1)))
        begin
          if ($unsigned(wire731))
            begin
              reg807 = ($signed((~reg440[(1'h1):(1'h0)])) ?
                  wire414[(2'h2):(2'h2)] : ((8'hba) ?
                      (~^reg798) : (forvar734 <= $signed(reg420[(1'h1):(1'h1)]))));
              reg808 <= (~|reg773);
              reg809 <= wire434[(2'h3):(2'h3)];
            end
          else
            begin
              reg807 <= ((($unsigned((reg739 >>> reg790)) == reg765) ?
                  ($unsigned({reg764}) ?
                      ((|forvar795) ?
                          $signed((8'hb6)) : $unsigned(reg740)) : $signed((forvar734 ?
                          wire416 : reg440))) : (&{forvar438[(2'h2):(1'h0)],
                      (~|wire413)})) | reg768[(2'h2):(2'h2)]);
              reg808 = (+reg800);
              reg809 <= "ELbmS4pipb1pDVuWams";
              reg810 = {($unsigned(reg736[(1'h1):(1'h0)]) * (((reg800 <= reg429) + (reg751 ?
                      forvar806 : wire418)) ^~ (7'h42)))};
            end
          reg811 <= reg792;
          for (forvar812 = (1'h0); (forvar812 < (2'h2)); forvar812 = (forvar812 + (1'h1)))
            begin
              reg813 <= $unsigned(($unsigned($unsigned($unsigned(reg421))) ~^ $signed((reg798[(3'h6):(3'h6)] + reg750))));
              reg814 = reg777;
              reg815 <= $unsigned((-$signed($unsigned($unsigned(reg783)))));
              reg816 <= $unsigned((&"mKQf5"));
            end
        end
      reg817 = wire731[(3'h5):(1'h1)];
      reg818 <= (reg762 ? reg784[(3'h4):(2'h3)] : $unsigned((7'h44)));
      for (forvar819 = (1'h0); (forvar819 < (3'h4)); forvar819 = (forvar819 + (1'h1)))
        begin
          for (forvar820 = (1'h0); (forvar820 < (2'h2)); forvar820 = (forvar820 + (1'h1)))
            begin
              reg821 = reg807;
              reg822 <= $unsigned($signed($unsigned($unsigned(forvar771))));
              reg823 <= $unsigned((forvar789[(4'hd):(2'h3)] ?
                  reg783 : ($unsigned({reg808, forvar789}) ?
                      wire416[(1'h1):(1'h1)] : {$unsigned(wire415)})));
              reg824 = (reg425 > (reg782[(2'h2):(2'h2)] ?
                  $signed(reg755) : $unsigned($unsigned("fZFBilg0"))));
            end
          if ($signed((reg748[(4'hf):(2'h2)] ?
              $unsigned((-(reg774 ?
                  wire441 : reg784))) : $unsigned(reg785[(1'h1):(1'h1)]))))
            begin
              reg825 <= $signed({$unsigned($unsigned((reg765 & forvar423)))});
            end
          else
            begin
              reg825 <= (-$unsigned((-{$unsigned(reg784),
                  (wire416 ? reg796 : (8'ha7))})));
              reg826 = ($signed((((|(8'hb8)) ? reg740 : (8'ha7)) ?
                      forvar799[(4'hb):(3'h5)] : reg763)) ?
                  ($unsigned((reg738[(5'h10):(3'h6)] ?
                      {reg439,
                          (8'haa)} : {reg780})) && reg736[(4'h8):(3'h4)]) : "5i2rCWG4k8epvtMW");
              reg827 <= ((((reg813[(1'h0):(1'h0)] || (|wire731)) + (8'hb7)) ?
                  "ITqbEGU" : ((8'hb0) | wire775)) < reg739[(3'h5):(3'h5)]);
            end
        end
    end
  assign wire828 = ((reg736[(3'h7):(2'h2)] < (((reg750 ?
                           reg748 : reg431) || (+reg773)) ?
                       {forvar422} : (((8'hbc) ? wire731 : reg772) ?
                           $unsigned(reg768) : (reg779 <<< reg773)))) > (reg827[(3'h6):(3'h6)] ?
                       ("RImNvIKyFC30LVH2Jsqm" ?
                           (^~(forvar758 ?
                               reg747 : (7'h43))) : reg419[(3'h6):(2'h3)]) : $unsigned((8'hab))));
  assign wire829 = $signed((reg431[(1'h1):(1'h0)] ?
                       (~^{$unsigned(reg809),
                           forvar819}) : $signed(((|(8'hbb)) ^~ wire416[(3'h6):(3'h4)]))));
  assign wire830 = ($unsigned((({forvar771,
                       reg428} >>> reg782) >> $unsigned(reg738))) * ((~reg737[(1'h0):(1'h0)]) ?
                       $signed($signed(reg769[(3'h7):(1'h0)])) : {reg787,
                           (8'haf)}));
  assign wire831 = ($signed(($signed($signed((8'hb3))) != $signed({wire830,
                           wire830}))) ?
                       (!reg740[(3'h5):(3'h4)]) : $unsigned(({(reg801 >> forvar789),
                               $signed(wire414)} ?
                           reg792 : ({reg737, wire416} ?
                               (reg755 ? reg439 : wire830) : reg803))));
  module832 modinst927 (.wire836(reg747), .wire833(reg769), .clk(clk), .y(wire926), .wire834(wire829), .wire835(reg825));
  assign wire928 = (reg784 | (~^$unsigned(($signed(reg801) && "5UcLb2hvB7FiSUD"))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module71
#( parameter param408 = ((((((8'hbb) == (8'h9c)) > (|(8'hbd))) ? (((8'ha3) ? (8'ha7) : (8'hbe)) > ((8'hab) << (8'hbf))) : (~|(8'ha9))) ? ((((8'hab) ? (8'hb0) : (8'had)) ? {(8'hab)} : ((8'hb4) | (8'ha0))) ? (&((8'had) ? (8'h9d) : (7'h44))) : {((8'h9e) ? (8'ha9) : (8'h9c)), (!(8'ha0))}) : (!((8'ha1) + (|(8'ha7))))) ? (8'ha0) : (({(8'hb6), {(7'h41)}} >>> (((8'ha2) ? (8'ha2) : (8'had)) ? {(8'hb4), (7'h40)} : {(8'hae)})) ? (8'ha1) : {(((8'ha9) << (8'ha2)) ? ((8'ha0) ? (8'hb0) : (8'ha0)) : ((8'hac) - (7'h44))), ({(8'hbd)} ^~ {(8'h9e), (8'hbf)})})) )
(y, clk, wire76, wire75, wire74, wire73, wire72);
  output wire [(32'h523):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire76;
  input wire [(2'h3):(1'h0)] wire75;
  input wire [(4'he):(1'h0)] wire74;
  input wire signed [(4'hd):(1'h0)] wire73;
  input wire signed [(4'hf):(1'h0)] wire72;
  wire signed [(4'ha):(1'h0)] wire407;
  wire [(4'ha):(1'h0)] wire406;
  wire [(4'h9):(1'h0)] wire405;
  reg signed [(5'h10):(1'h0)] reg400 = (1'h0);
  reg [(2'h2):(1'h0)] forvar395 = (1'h0);
  reg [(4'h9):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg404 = (1'h0);
  reg [(5'h13):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg402 = (1'h0);
  reg [(3'h7):(1'h0)] reg401 = (1'h0);
  reg [(4'hf):(1'h0)] forvar400 = (1'h0);
  reg [(2'h2):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg397 = (1'h0);
  reg [(5'h14):(1'h0)] reg396 = (1'h0);
  reg [(5'h11):(1'h0)] reg395 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg394 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar393 = (1'h0);
  reg [(3'h6):(1'h0)] reg392 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire391;
  wire signed [(3'h7):(1'h0)] wire264;
  wire signed [(4'hf):(1'h0)] wire140;
  reg [(4'h9):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg137 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg136 = (1'h0);
  reg [(5'h12):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar132 = (1'h0);
  reg [(5'h12):(1'h0)] reg131 = (1'h0);
  reg [(4'hc):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg129 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg128 = (1'h0);
  reg [(3'h7):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg126 = (1'h0);
  reg [(2'h3):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg124 = (1'h0);
  reg [(2'h2):(1'h0)] forvar123 = (1'h0);
  reg [(3'h7):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg121 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg118 = (1'h0);
  reg [(3'h4):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg116 = (1'h0);
  reg [(5'h15):(1'h0)] forvar115 = (1'h0);
  reg [(4'hd):(1'h0)] forvar114 = (1'h0);
  wire [(4'h9):(1'h0)] wire113;
  wire signed [(5'h15):(1'h0)] wire112;
  reg [(4'h8):(1'h0)] reg111 = (1'h0);
  reg [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg109 = (1'h0);
  reg [(3'h5):(1'h0)] reg108 = (1'h0);
  reg [(3'h5):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar106 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar105 = (1'h0);
  wire [(3'h4):(1'h0)] wire104;
  wire signed [(5'h12):(1'h0)] wire103;
  reg signed [(4'h8):(1'h0)] reg102 = (1'h0);
  reg [(5'h14):(1'h0)] reg101 = (1'h0);
  reg [(4'ha):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar99 = (1'h0);
  reg [(4'h8):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg97 = (1'h0);
  reg [(4'ha):(1'h0)] forvar96 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg95 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg94 = (1'h0);
  reg [(5'h10):(1'h0)] reg93 = (1'h0);
  reg [(4'hb):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar91 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg90 = (1'h0);
  reg [(3'h7):(1'h0)] reg89 = (1'h0);
  reg [(5'h13):(1'h0)] reg88 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar85 = (1'h0);
  reg [(3'h5):(1'h0)] reg84 = (1'h0);
  reg [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg82 = (1'h0);
  reg [(2'h3):(1'h0)] forvar81 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar79 = (1'h0);
  wire [(4'hf):(1'h0)] wire78;
  wire signed [(5'h14):(1'h0)] wire77;
  wire signed [(4'hf):(1'h0)] wire266;
  reg signed [(3'h4):(1'h0)] forvar267 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar269 = (1'h0);
  reg [(3'h5):(1'h0)] reg270 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg271 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg272 = (1'h0);
  reg [(3'h7):(1'h0)] reg273 = (1'h0);
  reg [(3'h6):(1'h0)] reg274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar276 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg277 = (1'h0);
  reg [(5'h14):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg279 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg280 = (1'h0);
  reg [(3'h5):(1'h0)] reg281 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg283 = (1'h0);
  reg [(4'hf):(1'h0)] reg284 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg285 = (1'h0);
  reg [(5'h10):(1'h0)] reg286 = (1'h0);
  reg [(4'h9):(1'h0)] reg287 = (1'h0);
  reg [(5'h15):(1'h0)] reg288 = (1'h0);
  reg [(5'h15):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg290 = (1'h0);
  reg [(5'h13):(1'h0)] reg291 = (1'h0);
  reg [(4'hc):(1'h0)] reg292 = (1'h0);
  reg [(5'h13):(1'h0)] reg293 = (1'h0);
  wire [(4'hb):(1'h0)] wire389;
  assign y = {wire407,
                 wire406,
                 wire405,
                 reg400,
                 forvar395,
                 reg393,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 forvar400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 reg392,
                 wire391,
                 wire264,
                 wire140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 forvar132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 forvar123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 forvar115,
                 forvar114,
                 wire113,
                 wire112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 forvar106,
                 forvar105,
                 wire104,
                 wire103,
                 reg102,
                 reg101,
                 reg100,
                 forvar99,
                 reg98,
                 reg97,
                 forvar96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 forvar91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 forvar85,
                 reg84,
                 reg83,
                 reg82,
                 forvar81,
                 reg80,
                 forvar79,
                 wire78,
                 wire77,
                 wire266,
                 forvar267,
                 reg268,
                 forvar269,
                 reg270,
                 reg271,
                 reg272,
                 reg273,
                 reg274,
                 reg275,
                 forvar276,
                 reg277,
                 reg278,
                 reg279,
                 reg280,
                 reg281,
                 forvar282,
                 reg283,
                 reg284,
                 reg285,
                 reg286,
                 reg287,
                 reg288,
                 reg289,
                 reg290,
                 reg291,
                 reg292,
                 reg293,
                 wire389,
                 (1'h0)};
  assign wire77 = $signed($unsigned(wire76[(1'h0):(1'h0)]));
  assign wire78 = wire74;
  always
    @(posedge clk) begin
      for (forvar79 = (1'h0); (forvar79 < (2'h3)); forvar79 = (forvar79 + (1'h1)))
        begin
          reg80 = $unsigned((~$signed($unsigned($signed(wire76)))));
          for (forvar81 = (1'h0); (forvar81 < (2'h3)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 <= wire77[(5'h11):(2'h3)];
              reg83 <= {reg80[(1'h1):(1'h0)]};
              reg84 = (((wire74[(4'h9):(2'h3)] && wire73[(4'h9):(4'h8)]) ?
                      wire75[(2'h2):(1'h1)] : (+wire78[(2'h3):(1'h0)])) ?
                  $unsigned(wire73[(4'hd):(3'h7)]) : reg80);
            end
        end
      for (forvar85 = (1'h0); (forvar85 < (1'h0)); forvar85 = (forvar85 + (1'h1)))
        begin
          if ({(~&(+(|forvar85))), (|$unsigned({(~^wire77)}))})
            begin
              reg86 <= reg83;
              reg87 <= $unsigned(wire74);
              reg88 = wire72[(2'h2):(1'h1)];
              reg89 = $unsigned(($signed($unsigned($unsigned(reg86))) ?
                  $signed(($unsigned((8'hab)) << reg82)) : reg80));
              reg90 <= $unsigned(($signed(($signed(reg80) >> (wire72 >>> wire78))) || reg86[(1'h0):(1'h0)]));
            end
          else
            begin
              reg86 <= {((reg88[(1'h1):(1'h1)] | wire72[(3'h6):(3'h5)]) << ({$unsigned(reg90)} > ($signed((8'ha2)) == (reg80 << reg82))))};
            end
          for (forvar91 = (1'h0); (forvar91 < (2'h2)); forvar91 = (forvar91 + (1'h1)))
            begin
              reg92 = ($signed($unsigned((~|forvar79))) ^~ forvar81[(2'h3):(2'h2)]);
            end
          reg93 <= (^~{(reg80 ? (~^((8'ha7) & reg90)) : $signed((^wire73))),
              ("sz8e" ? reg86[(1'h1):(1'h1)] : {$unsigned(forvar81)})});
        end
      reg94 <= wire72[(2'h2):(1'h1)];
      reg95 = $signed(reg84[(1'h0):(1'h0)]);
      for (forvar96 = (1'h0); (forvar96 < (1'h1)); forvar96 = (forvar96 + (1'h1)))
        begin
          reg97 <= reg84;
          reg98 <= (+forvar91);
          for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 = (~(!(~^$signed($unsigned(reg95)))));
              reg101 = (wire74 ^~ ($unsigned(({(8'ha2),
                      reg89} > $signed(wire73))) ?
                  ({$signed(reg97), wire74} ?
                      reg80 : ({reg86} != (reg100 ?
                          forvar99 : reg82))) : $unsigned((!forvar79))));
            end
          reg102 = (~&wire76[(3'h4):(1'h0)]);
        end
    end
  assign wire103 = (!(wire75[(1'h0):(1'h0)] ? "Ri" : reg88[(3'h4):(1'h1)]));
  assign wire104 = (~^(~|forvar81[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar105 = (1'h0); (forvar105 < (3'h4)); forvar105 = (forvar105 + (1'h1)))
        begin
          for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 <= (8'ha4);
            end
          reg108 <= {$signed((~|$signed((reg86 ? reg82 : wire74))))};
          reg109 = $signed(wire104[(2'h2):(1'h0)]);
          reg110 <= (&reg100);
        end
      reg111 <= $unsigned(forvar81);
    end
  assign wire112 = (!forvar81[(2'h2):(2'h2)]);
  assign wire113 = (reg82[(4'hb):(1'h1)] - reg107[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar114 = (1'h0); (forvar114 < (2'h3)); forvar114 = (forvar114 + (1'h1)))
        begin
          for (forvar115 = (1'h0); (forvar115 < (2'h3)); forvar115 = (forvar115 + (1'h1)))
            begin
              reg116 = reg97;
              reg117 <= (-(^((7'h40) ?
                  {((7'h44) ? reg94 : (8'hbc)),
                      (-wire103)} : (!(reg97 + reg102)))));
              reg118 <= {((((forvar81 << reg102) ?
                          {forvar106, (8'h9c)} : (~^reg84)) ?
                      (~"pCYhQLoiA") : $unsigned(reg87[(1'h1):(1'h0)])) ~^ $signed(wire78[(4'hd):(3'h6)]))};
            end
          if (reg95[(3'h4):(1'h1)])
            begin
              reg119 = (&wire73);
            end
          else
            begin
              reg119 <= reg86;
              reg120 = reg101[(2'h3):(2'h2)];
              reg121 = (reg108[(2'h3):(2'h3)] >= {$signed((reg95[(1'h0):(1'h0)] * {wire113}))});
              reg122 = $signed({reg118});
            end
          for (forvar123 = (1'h0); (forvar123 < (1'h0)); forvar123 = (forvar123 + (1'h1)))
            begin
              reg124 = forvar79;
              reg125 = $unsigned({$unsigned(($unsigned(reg124) ?
                      (reg116 | reg117) : (reg118 ? reg101 : (7'h41)))),
                  wire74[(3'h6):(3'h5)]});
              reg126 = ({(wire77 ?
                      (|(forvar106 ?
                          reg87 : (7'h40))) : forvar114[(2'h2):(1'h0)]),
                  $unsigned({(~^reg89),
                      (~^wire103)})} >>> reg87[(1'h0):(1'h0)]);
              reg127 <= ((($unsigned((reg94 ?
                          reg119 : (8'hac))) >>> $signed({reg119, wire112})) ?
                      $unsigned("5pFm2Wb8w3gYhsB") : (-forvar123)) ?
                  (~^reg94[(1'h1):(1'h1)]) : (+$unsigned(((~(8'ha5)) >> ((8'hbb) ?
                      (8'ha0) : wire75)))));
            end
        end
      if ($unsigned({(reg116 & (reg125[(1'h1):(1'h1)] ?
              (reg117 | reg84) : (forvar105 ? reg98 : (8'hb3)))),
          $signed(wire113)}))
        begin
          if ((~^(&(+reg90[(1'h0):(1'h0)]))))
            begin
              reg128 = reg95[(3'h4):(3'h4)];
              reg129 = ((-(forvar99 & $unsigned((wire113 && wire104)))) <= reg108);
              reg130 = $signed(reg101);
            end
          else
            begin
              reg128 <= "zgBbvkBVREg";
              reg129 = reg126[(4'he):(4'he)];
              reg130 = (~|wire78);
              reg131 <= $unsigned($signed((~^(^~(reg101 ? wire78 : reg117)))));
            end
          for (forvar132 = (1'h0); (forvar132 < (1'h1)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 = reg92;
              reg134 <= {reg98};
              reg135 <= (~|(8'hb2));
              reg136 = reg108[(1'h0):(1'h0)];
              reg137 <= {$unsigned($unsigned(("O9qfbLYds4dGFRrdAxDw" | reg101[(2'h2):(1'h1)]))),
                  $signed($unsigned((forvar79 ?
                      reg82[(4'hc):(3'h6)] : $unsigned(reg128))))};
            end
          reg138 = "pWfw6Ecdsatb8X2";
          reg139 = $signed((8'hbf));
        end
      else
        begin
          if (reg119[(1'h0):(1'h0)])
            begin
              reg128 <= (($signed(($unsigned(forvar115) & (forvar105 * forvar81))) ?
                      reg128[(4'hb):(3'h4)] : $signed((^~reg119[(3'h7):(1'h1)]))) ?
                  (+reg87) : ((^~$unsigned({forvar91})) ?
                      (&(|(8'hba))) : reg128));
              reg129 <= reg86[(1'h0):(1'h0)];
              reg130 = ((((+$unsigned(reg129)) ?
                          forvar81[(2'h2):(2'h2)] : {(|reg89)}) ?
                      reg82[(4'he):(3'h7)] : (~|(~(^~reg87)))) ?
                  reg137[(5'h14):(4'hc)] : "Ww");
              reg131 = {reg117[(2'h3):(1'h0)], reg138[(3'h6):(2'h3)]};
            end
          else
            begin
              reg128 = reg133[(3'h7):(1'h1)];
              reg129 = $signed((reg97 >>> {((8'hb1) <= {reg109}),
                  $signed({reg89})}));
              reg130 <= ($unsigned((reg93 ?
                      reg119[(4'hc):(2'h3)] : $unsigned($unsigned(reg136)))) ?
                  $unsigned($unsigned((~|{wire74}))) : wire73[(3'h6):(1'h0)]);
            end
          for (forvar132 = (1'h0); (forvar132 < (3'h4)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= reg120[(2'h2):(2'h2)];
            end
          reg134 <= ({(|((wire74 || reg138) ?
                      $signed(reg97) : (reg93 - (7'h42))))} ?
              (((8'hb4) ?
                      $signed(reg126[(4'hb):(2'h2)]) : reg86[(1'h1):(1'h0)]) ?
                  (($unsigned(reg110) - {(8'ha9)}) - {(~&(8'haf))}) : ("xkAP" | "S9m0GX1QTVNbK65NKU0g")) : $signed(reg107));
          reg135 = $signed($signed(wire104[(3'h4):(2'h3)]));
          reg136 = reg88;
        end
    end
  assign wire140 = (~wire75);
  module141 modinst265 (wire264, clk, forvar79, reg93, reg137, reg109, forvar91);
  assign wire266 = (!reg90[(4'hb):(1'h0)]);
  always
    @(posedge clk) begin
      for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
        begin
          reg268 = $unsigned($unsigned($unsigned(($unsigned(reg119) ?
              wire73 : reg90))));
        end
      for (forvar269 = (1'h0); (forvar269 < (2'h2)); forvar269 = (forvar269 + (1'h1)))
        begin
          reg270 = $signed((&{($unsigned((8'hb9)) ?
                  $signed((7'h44)) : (|wire264)),
              {(reg137 ? wire266 : (7'h43)), reg95[(2'h3):(1'h0)]}}));
        end
      if ($unsigned(reg139))
        begin
          reg271 <= {reg108[(1'h1):(1'h1)]};
        end
      else
        begin
          if (reg83)
            begin
              reg271 = (&forvar123);
              reg272 <= {($unsigned({(reg138 != reg87)}) == ($unsigned(reg136) ?
                      ((|reg139) ?
                          {reg110,
                              reg130} : ((7'h40) ~^ forvar267)) : (reg133[(2'h2):(1'h1)] ?
                          (^~reg129) : $unsigned(forvar81)))),
                  $unsigned((~&$signed(reg110[(3'h5):(1'h0)])))};
              reg273 = ($unsigned((~&$signed(forvar81))) ?
                  (~^$unsigned(forvar106[(4'hd):(4'hc)])) : reg109);
              reg274 = {$unsigned(reg107[(3'h4):(1'h0)])};
            end
          else
            begin
              reg271 = $unsigned({$unsigned(forvar99[(3'h6):(2'h2)]),
                  $signed((((7'h43) ? reg107 : reg139) != $signed(reg134)))});
              reg272 <= (~^$signed((~|(~&$unsigned(forvar91)))));
            end
          reg275 <= ($signed((wire104[(2'h2):(2'h2)] >> ("W5oVA4dvPbyvG8" ?
              $signed(reg108) : ((8'hba) ? (8'hb9) : (8'hbd))))) != (~(8'hbc)));
          for (forvar276 = (1'h0); (forvar276 < (2'h3)); forvar276 = (forvar276 + (1'h1)))
            begin
              reg277 <= {(reg82 ?
                      ({(forvar91 ? forvar132 : reg109), "VDeUZtkT5"} ?
                          {{reg107, forvar96},
                              (reg94 ^~ forvar96)} : (|(reg133 ^~ (8'hb0)))) : (((reg117 ?
                              reg110 : forvar123) >> reg273[(3'h6):(1'h1)]) ?
                          reg135 : (~$unsigned(forvar91)))),
                  reg107[(1'h0):(1'h0)]};
              reg278 <= (!$unsigned(reg80[(1'h1):(1'h1)]));
              reg279 <= ($signed({$signed(reg130)}) >> ((~((|(8'ha5)) >= (forvar106 < reg270))) < (-($signed((8'hb2)) ?
                  $unsigned((8'hac)) : reg84))));
              reg280 = forvar132;
              reg281 = $signed((+(({(8'haa),
                  forvar91} ^~ wire74) >= ((|reg279) ?
                  $signed((8'haa)) : (reg272 ^~ reg125)))));
            end
          for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
            begin
              reg283 <= (-reg279[(1'h1):(1'h0)]);
              reg284 = reg134;
              reg285 <= ($unsigned($signed($unsigned((reg128 ?
                  (8'hba) : wire264)))) ^ $signed({($signed(reg124) ?
                      reg118[(1'h1):(1'h1)] : $signed(reg117)),
                  reg139}));
              reg286 <= (((!$signed($unsigned(forvar123))) ?
                  reg100[(4'h9):(1'h1)] : $unsigned({(reg284 && wire264)})) >= $signed($signed((&wire72))));
              reg287 <= reg275[(4'hc):(2'h3)];
            end
          reg288 = (-($signed(((reg84 ?
                  reg117 : wire140) ^ $unsigned(reg133))) ?
              {{$unsigned(reg83), $signed(wire72)}} : (reg120 ?
                  reg86 : {(reg128 <= reg135)})));
        end
    end
  always
    @(posedge clk) begin
      reg289 = reg268;
      reg290 <= $unsigned((^~(reg139 < ($signed(reg94) ?
          (-reg90) : ((8'hb3) ? (8'h9c) : reg131)))));
      reg291 = reg93;
      reg292 = (~^$unsigned($signed($signed(reg109[(1'h1):(1'h1)]))));
      reg293 = ($unsigned(reg131) || $unsigned({(~|reg127)}));
    end
  module294 modinst390 (.wire296(wire75), .wire298(wire73), .clk(clk), .wire299(reg137), .wire295(reg101), .y(wire389), .wire297(wire266));
  assign wire391 = $signed((($signed({(8'ha8)}) ?
                       (8'h9e) : wire266[(4'hd):(1'h1)]) + $signed((8'hb3))));
  always
    @(posedge clk) begin
      if ($unsigned({reg136[(1'h0):(1'h0)], reg138[(4'h9):(1'h0)]}))
        begin
          reg392 <= (-reg120[(1'h1):(1'h0)]);
          for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= reg130;
              reg395 = (^(reg87 ?
                  reg109[(4'hc):(2'h3)] : ($signed(wire391[(3'h7):(2'h2)]) ?
                      "H" : $unsigned(reg288[(5'h12):(4'h9)]))));
              reg396 <= reg119[(3'h4):(1'h0)];
              reg397 = (reg134 >>> reg290[(3'h4):(1'h1)]);
              reg398 = $signed($unsigned($unsigned(reg120[(1'h1):(1'h1)])));
            end
          reg399 = "QPleNARwp6KkCaoBa";
          for (forvar400 = (1'h0); (forvar400 < (2'h3)); forvar400 = (forvar400 + (1'h1)))
            begin
              reg401 = (~|$signed((+$unsigned(reg280[(1'h1):(1'h0)]))));
              reg402 <= ($signed(($signed((wire140 >>> reg394)) ?
                      $signed((forvar91 ? reg129 : forvar276)) : (8'h9d))) ?
                  {(forvar269[(4'ha):(2'h2)] ?
                          "ZLkYy" : (((8'hbb) ? reg88 : reg102) ?
                              $signed(forvar267) : (reg401 || reg286))),
                      $signed(((reg117 ? reg120 : reg289) ?
                          (!reg288) : (~^reg88)))} : (wire104 - wire74[(1'h0):(1'h0)]));
              reg403 <= reg95;
              reg404 <= $unsigned(reg92);
            end
        end
      else
        begin
          if ($unsigned(reg287))
            begin
              reg392 <= $unsigned(((reg392[(3'h5):(3'h5)] ?
                      reg394 : (!$unsigned(wire140))) ?
                  reg271 : $unsigned(reg95[(2'h2):(1'h0)])));
              reg393 <= (&(reg107 <<< $signed(((!reg110) ?
                  reg126[(4'he):(2'h3)] : wire104[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg392 <= ((7'h41) ?
                  (reg92[(3'h4):(3'h4)] ?
                      (wire103[(3'h5):(1'h0)] ~^ {((8'hab) | wire113)}) : $unsigned(reg392)) : wire266);
              reg393 = "Z8WJx8iqruxedK";
              reg394 <= "b7hfl8V81INusHS0C";
            end
          for (forvar395 = (1'h0); (forvar395 < (2'h2)); forvar395 = (forvar395 + (1'h1)))
            begin
              reg396 = $signed((!{$signed((reg82 >>> reg130)),
                  $unsigned((reg108 ? (8'h9c) : reg283))}));
            end
          if ((reg126 ? reg403 : (7'h42)))
            begin
              reg397 <= (8'hb1);
              reg398 = {(^~reg127),
                  (~&$signed(({forvar395, reg102} ?
                      reg392[(3'h6):(2'h2)] : {reg404, (8'hbf)})))};
              reg399 = reg80;
              reg400 = $signed(reg88);
            end
          else
            begin
              reg397 <= (!reg402[(1'h0):(1'h0)]);
              reg398 = reg93;
              reg399 <= "hziP7U94z4";
              reg400 = {((8'hbf) * {(|(^~(8'hac))), (~&reg95)})};
              reg401 = $unsigned((&reg124));
            end
        end
    end
  assign wire405 = $signed($unsigned({$signed(reg98)}));
  assign wire406 = (-{reg291[(5'h12):(3'h4)], (8'h9c)});
  assign wire407 = (reg101[(3'h7):(1'h0)] - $signed((reg128[(4'hb):(4'h8)] & (7'h40))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module294
#( parameter param387 = ((((~(8'hb0)) ? {((8'hb5) ~^ (8'h9f))} : (~^((8'ha7) < (8'haf)))) || ({((8'ha4) ? (8'ha4) : (8'hbb)), (^(8'haa))} == (|((8'haa) ? (8'ha0) : (8'ha9))))) < (|(~&(|(|(8'ha2))))))
, parameter param388 = param387 )
(y, clk, wire299, wire298, wire297, wire296, wire295);
  output wire [(32'h42b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire299;
  input wire [(3'h4):(1'h0)] wire298;
  input wire signed [(3'h4):(1'h0)] wire297;
  input wire [(2'h2):(1'h0)] wire296;
  input wire signed [(5'h14):(1'h0)] wire295;
  reg [(3'h5):(1'h0)] reg386 = (1'h0);
  reg [(4'hb):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg384 = (1'h0);
  reg [(4'ha):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar375 = (1'h0);
  reg [(3'h7):(1'h0)] reg383 = (1'h0);
  reg [(4'h8):(1'h0)] forvar382 = (1'h0);
  reg [(5'h14):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg380 = (1'h0);
  reg [(4'h8):(1'h0)] reg379 = (1'h0);
  reg [(2'h2):(1'h0)] reg378 = (1'h0);
  reg [(5'h13):(1'h0)] reg377 = (1'h0);
  reg [(5'h11):(1'h0)] reg376 = (1'h0);
  reg [(3'h7):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg374 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire373;
  wire [(5'h10):(1'h0)] wire372;
  wire [(4'hf):(1'h0)] wire371;
  wire [(4'h8):(1'h0)] wire370;
  reg signed [(4'hd):(1'h0)] reg369 = (1'h0);
  reg [(3'h5):(1'h0)] reg368 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire367;
  wire [(5'h12):(1'h0)] wire366;
  wire [(3'h6):(1'h0)] wire365;
  reg signed [(4'h8):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg362 = (1'h0);
  reg [(4'ha):(1'h0)] forvar361 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar360 = (1'h0);
  reg [(5'h13):(1'h0)] reg359 = (1'h0);
  reg [(3'h6):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg356 = (1'h0);
  reg [(5'h10):(1'h0)] forvar355 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg354 = (1'h0);
  reg [(4'hc):(1'h0)] reg353 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire352;
  reg [(5'h12):(1'h0)] reg351 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg350 = (1'h0);
  reg [(4'hc):(1'h0)] reg349 = (1'h0);
  reg signed [(4'he):(1'h0)] reg348 = (1'h0);
  reg [(5'h12):(1'h0)] forvar347 = (1'h0);
  reg [(2'h3):(1'h0)] reg346 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar345 = (1'h0);
  reg [(2'h3):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg343 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire342;
  reg [(4'h9):(1'h0)] reg341 = (1'h0);
  reg [(5'h13):(1'h0)] reg340 = (1'h0);
  reg [(3'h4):(1'h0)] reg339 = (1'h0);
  reg [(5'h11):(1'h0)] reg338 = (1'h0);
  reg [(2'h3):(1'h0)] forvar337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg336 = (1'h0);
  reg [(3'h5):(1'h0)] reg335 = (1'h0);
  reg [(3'h4):(1'h0)] forvar330 = (1'h0);
  reg [(4'hf):(1'h0)] forvar327 = (1'h0);
  reg [(4'hd):(1'h0)] reg334 = (1'h0);
  reg [(5'h13):(1'h0)] reg333 = (1'h0);
  reg [(4'he):(1'h0)] reg332 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg331 = (1'h0);
  reg [(2'h3):(1'h0)] reg330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg329 = (1'h0);
  reg [(5'h13):(1'h0)] reg328 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg327 = (1'h0);
  reg [(3'h5):(1'h0)] reg326 = (1'h0);
  reg [(4'hd):(1'h0)] reg325 = (1'h0);
  reg [(4'hb):(1'h0)] reg324 = (1'h0);
  reg [(4'hd):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg321 = (1'h0);
  reg [(4'h9):(1'h0)] forvar320 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg319 = (1'h0);
  reg [(3'h6):(1'h0)] forvar318 = (1'h0);
  reg [(4'hd):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg316 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg315 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar314 = (1'h0);
  reg [(5'h14):(1'h0)] reg312 = (1'h0);
  reg [(5'h15):(1'h0)] reg313 = (1'h0);
  reg [(5'h12):(1'h0)] forvar312 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg311 = (1'h0);
  reg [(5'h14):(1'h0)] reg310 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar309 = (1'h0);
  reg [(3'h6):(1'h0)] reg308 = (1'h0);
  reg [(4'hb):(1'h0)] reg307 = (1'h0);
  reg [(3'h6):(1'h0)] reg306 = (1'h0);
  reg [(2'h3):(1'h0)] reg305 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg304 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg303 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire302;
  wire [(4'h9):(1'h0)] wire301;
  wire [(5'h10):(1'h0)] wire300;
  assign y = {reg386,
                 reg385,
                 reg384,
                 reg382,
                 forvar375,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 wire373,
                 wire372,
                 wire371,
                 wire370,
                 reg369,
                 reg368,
                 wire367,
                 wire366,
                 wire365,
                 reg364,
                 reg363,
                 reg362,
                 forvar361,
                 forvar360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 forvar355,
                 reg354,
                 reg353,
                 wire352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 forvar347,
                 reg346,
                 forvar345,
                 reg344,
                 reg343,
                 wire342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 forvar337,
                 reg336,
                 reg335,
                 forvar330,
                 forvar327,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 forvar318,
                 reg317,
                 reg316,
                 reg315,
                 forvar314,
                 reg312,
                 reg313,
                 forvar312,
                 reg311,
                 reg310,
                 forvar309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 wire302,
                 wire301,
                 wire300,
                 (1'h0)};
  assign wire300 = wire297;
  assign wire301 = $unsigned(wire296[(1'h1):(1'h0)]);
  assign wire302 = $unsigned((|wire301[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      reg303 <= ({(wire301 ~^ "YoiCpFs6BWNCgo6")} && $unsigned(wire295));
      if (($signed($signed(wire297[(1'h0):(1'h0)])) ?
          wire302[(3'h7):(3'h5)] : wire300[(4'hd):(2'h2)]))
        begin
          if ((wire302 != wire300))
            begin
              reg304 <= {$unsigned($signed((!(wire298 - wire298)))),
                  {"Owtkmn8LdutIOf"}};
              reg305 <= wire296;
              reg306 = (($signed({wire300[(2'h2):(1'h0)], $signed(reg305)}) ?
                  ("AlSvcQdwDZ2hOuRGECQL" ?
                      (&(wire295 ?
                          reg304 : (8'had))) : $signed($signed(wire302))) : reg305[(2'h3):(1'h1)]) != $signed((wire298 ?
                  $signed(wire296) : $signed((8'hab)))));
              reg307 = $unsigned((wire302[(3'h4):(2'h3)] != reg306));
              reg308 = $signed("kBQiIqpMXaCX");
            end
          else
            begin
              reg304 <= {wire296};
              reg305 <= {((({wire298} ?
                      (reg303 * (8'hbd)) : (reg307 ?
                          wire297 : reg305)) >> wire295) * $signed("")),
                  {reg303[(2'h3):(1'h1)]}};
            end
          for (forvar309 = (1'h0); (forvar309 < (1'h0)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 = wire300[(3'h6):(3'h5)];
              reg311 <= (!reg308);
            end
          for (forvar312 = (1'h0); (forvar312 < (3'h4)); forvar312 = (forvar312 + (1'h1)))
            begin
              reg313 = {forvar309[(1'h1):(1'h1)]};
            end
        end
      else
        begin
          if ((-reg304))
            begin
              reg304 <= $signed((~|({(wire295 ?
                      wire301 : (8'h9c))} << forvar312[(4'ha):(4'h8)])));
              reg305 = ((-{forvar312, {(^~reg307)}}) & wire295[(3'h4):(2'h3)]);
              reg306 <= $signed((+($signed((wire301 ? (8'ha9) : wire298)) ?
                  (~^(wire301 ? wire298 : reg311)) : $unsigned(((8'had) ?
                      reg304 : (8'ha2))))));
              reg307 <= (-(($signed($unsigned((7'h42))) | reg303[(2'h2):(2'h2)]) - {(((8'hba) ?
                      (8'haf) : forvar312) * reg310)}));
              reg308 = (^~reg310);
            end
          else
            begin
              reg304 <= wire295[(5'h12):(4'hb)];
            end
          for (forvar309 = (1'h0); (forvar309 < (2'h3)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 = (&$unsigned((reg303[(1'h0):(1'h0)] ?
                  ({wire302, forvar309} > $signed((7'h43))) : (~^(wire299 ?
                      reg313 : (8'hbd))))));
            end
          reg311 <= $signed(reg311[(2'h3):(2'h3)]);
          if (reg308[(1'h0):(1'h0)])
            begin
              reg312 = reg303;
              reg313 <= $signed({forvar309});
            end
          else
            begin
              reg312 = wire299[(3'h7):(3'h4)];
              reg313 = reg308[(2'h2):(1'h1)];
            end
          for (forvar314 = (1'h0); (forvar314 < (2'h3)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg315 = (wire299 ? reg305 : ({"Gx8YINQpZJczQkpT"} >> wire300));
              reg316 = $signed("pXURCt");
              reg317 = reg303[(1'h1):(1'h1)];
            end
        end
      for (forvar318 = (1'h0); (forvar318 < (2'h3)); forvar318 = (forvar318 + (1'h1)))
        begin
          reg319 <= (~(~&((8'ha4) + wire296)));
          for (forvar320 = (1'h0); (forvar320 < (1'h0)); forvar320 = (forvar320 + (1'h1)))
            begin
              reg321 <= (wire302 ^ {$unsigned($signed((~|wire297))),
                  $signed({forvar312})});
              reg322 = {reg311, "qXOq2LMVH"};
              reg323 <= (-reg311[(1'h1):(1'h0)]);
              reg324 <= $unsigned((&$signed($signed((wire296 ?
                  (8'hbe) : reg312)))));
            end
        end
      reg325 <= $unsigned(reg306);
    end
  always
    @(posedge clk) begin
      if (reg319[(1'h0):(1'h0)])
        begin
          reg326 <= reg304;
          if (wire302[(4'h9):(3'h4)])
            begin
              reg327 <= $signed(((reg308[(3'h5):(2'h2)] >> reg322) << $unsigned(("0rTG3nVBDG7HMe" >= $signed((8'h9f))))));
            end
          else
            begin
              reg327 = $signed(forvar318[(3'h4):(2'h3)]);
            end
          if ((^~wire302))
            begin
              reg328 <= wire295[(1'h0):(1'h0)];
              reg329 <= reg304[(2'h3):(1'h0)];
              reg330 = reg323[(2'h2):(1'h0)];
            end
          else
            begin
              reg328 = (^~$unsigned(reg324[(1'h0):(1'h0)]));
              reg329 = (~&(~^$unsigned("S1")));
              reg330 = (($signed($unsigned("rNzhc0bnSJA8ZDXXvG")) ^~ ($unsigned(forvar309[(4'ha):(4'ha)]) ?
                      $signed((~reg321)) : $unsigned($signed(reg321)))) ?
                  $unsigned($unsigned(({forvar314,
                      (8'h9f)} << $signed(wire297)))) : {(($signed(forvar312) & $unsigned(reg315)) > (reg305 < reg327[(3'h4):(2'h2)]))});
            end
          if ({(($signed({reg328}) == ((+(8'h9c)) ?
                  ((8'h9f) ? reg328 : forvar309) : (&reg319))) >= reg317),
              (8'ha6)})
            begin
              reg331 = reg316[(3'h7):(2'h2)];
            end
          else
            begin
              reg331 <= wire299;
              reg332 <= (forvar320[(3'h7):(3'h6)] ?
                  ((reg328 ?
                          reg324 : ((wire302 > reg308) >> (reg311 ~^ reg310))) ?
                      $signed($signed($signed(reg312))) : (((reg326 ?
                          reg329 : reg326) ^ $unsigned(wire295)) >> ($unsigned(reg310) ?
                          (forvar314 ?
                              wire302 : reg305) : forvar309[(4'hb):(4'ha)]))) : ("da" ?
                      wire297[(3'h4):(1'h0)] : ((forvar312[(4'h8):(2'h3)] <= $signed(forvar314)) ?
                          $unsigned((+reg311)) : (~^(reg325 << forvar314)))));
              reg333 <= ((wire299 ?
                      wire301[(4'h9):(3'h4)] : {((reg329 >>> forvar318) ?
                              "zdPeaMlaUXBsGIrac1" : reg317[(3'h5):(2'h2)])}) ?
                  reg322[(4'h8):(4'h8)] : ((reg324 < $unsigned((reg322 && wire302))) ?
                      (reg332[(3'h7):(1'h1)] ?
                          (reg328[(4'h9):(1'h0)] || (forvar312 << reg317)) : ($unsigned(reg317) ?
                              forvar320 : (reg321 >= reg315))) : ((~|(reg331 ?
                          reg308 : (8'ha2))) <= (8'hab))));
              reg334 = $unsigned((reg304[(2'h2):(2'h2)] >> $unsigned(reg327[(2'h2):(2'h2)])));
            end
        end
      else
        begin
          reg326 = reg311;
          for (forvar327 = (1'h0); (forvar327 < (2'h2)); forvar327 = (forvar327 + (1'h1)))
            begin
              reg328 <= forvar314;
              reg329 <= (&wire295[(1'h0):(1'h0)]);
            end
          for (forvar330 = (1'h0); (forvar330 < (1'h0)); forvar330 = (forvar330 + (1'h1)))
            begin
              reg331 <= ($signed(forvar330) ?
                  "Wpg9CLCbdA8QkW" : $unsigned(($unsigned($signed(reg303)) >> forvar314[(4'h8):(1'h0)])));
              reg332 <= $unsigned(reg307[(3'h6):(2'h2)]);
              reg333 = "hYP";
            end
        end
      if ($signed(((^~forvar320[(3'h4):(3'h4)]) ?
          (($signed((8'hbb)) ? {reg308, reg327} : ((8'haa) * reg334)) ?
              ($signed((8'hb4)) ?
                  (wire300 + reg303) : {reg322}) : $unsigned($signed(reg316))) : {($unsigned(reg325) ?
                  $unsigned(forvar314) : {wire302})})))
        begin
          reg335 <= (+reg312[(5'h14):(2'h2)]);
        end
      else
        begin
          reg335 <= reg332;
          reg336 <= ((|forvar314[(1'h1):(1'h1)]) & {(^~wire298[(2'h3):(1'h1)])});
          for (forvar337 = (1'h0); (forvar337 < (1'h1)); forvar337 = (forvar337 + (1'h1)))
            begin
              reg338 <= (({{(wire295 ^~ forvar320), {(8'hb8)}}} ?
                      reg322 : $signed((8'hbe))) ?
                  {{reg334[(3'h6):(3'h5)],
                          ((8'hb1) & (forvar320 ? reg336 : reg310))},
                      {$unsigned(reg331),
                          (!(forvar320 <<< forvar309))}} : (-$unsigned($unsigned((reg334 * wire295)))));
              reg339 = $unsigned($signed(wire300[(4'he):(3'h4)]));
              reg340 <= reg321;
              reg341 <= $signed("dpPLD15");
            end
        end
    end
  assign wire342 = $unsigned($signed((reg304[(2'h3):(1'h1)] << reg313[(3'h4):(1'h0)])));
  always
    @(posedge clk) begin
      reg343 <= forvar337;
      reg344 <= ((&(~|forvar330)) ?
          $signed(reg330[(2'h2):(2'h2)]) : reg307[(2'h2):(1'h0)]);
      for (forvar345 = (1'h0); (forvar345 < (1'h1)); forvar345 = (forvar345 + (1'h1)))
        begin
          reg346 = (reg321[(1'h0):(1'h0)] + $unsigned(wire298));
          for (forvar347 = (1'h0); (forvar347 < (1'h0)); forvar347 = (forvar347 + (1'h1)))
            begin
              reg348 = reg324;
              reg349 = reg328;
              reg350 <= ((~(~{$signed((8'hbd)), reg328[(4'hf):(4'hc)]})) ?
                  $signed(reg344[(1'h1):(1'h1)]) : ((&wire342) ?
                      (~^{((8'hb9) ~^ reg334)}) : (reg344[(1'h0):(1'h0)] ?
                          "oFqp" : $unsigned((reg303 ? reg344 : reg341)))));
            end
        end
      reg351 <= ($signed(($signed(reg339) >= ((-reg322) ?
              forvar314 : (!reg326)))) ?
          $unsigned((-reg312[(5'h13):(4'h9)])) : $unsigned(reg324[(4'h9):(3'h7)]));
    end
  assign wire352 = $signed((^(wire299[(4'h8):(1'h1)] >>> $signed(reg330))));
  always
    @(posedge clk) begin
      reg353 <= ($unsigned($signed(($signed(reg319) ?
              (reg316 > reg328) : (reg329 < reg310)))) ?
          (&$signed(((^reg350) & (forvar347 <= reg338)))) : (wire342 ?
              {(~&(forvar330 ^ reg349))} : reg340));
      reg354 <= (reg310 <= (reg303[(2'h2):(1'h0)] ?
          {reg311[(1'h0):(1'h0)]} : {((~^reg316) ^~ reg319[(3'h5):(3'h5)])}));
      for (forvar355 = (1'h0); (forvar355 < (1'h0)); forvar355 = (forvar355 + (1'h1)))
        begin
          reg356 <= $unsigned(((~|reg306[(3'h5):(2'h2)]) | reg303));
        end
      if ($signed(wire302))
        begin
          reg357 <= ($signed((8'hba)) & (+(^reg304[(3'h6):(2'h2)])));
          reg358 = ($unsigned((reg307 >>> ($unsigned(reg346) >> reg339[(2'h3):(2'h3)]))) * (((~((8'h9f) > reg340)) ?
              $signed(reg322[(5'h10):(4'ha)]) : forvar327) <<< (&$unsigned((!reg353)))));
          reg359 <= reg350[(4'h9):(3'h5)];
        end
      else
        begin
          reg357 = ({((forvar309[(1'h0):(1'h0)] >> {reg359, reg353}) ?
                      forvar330 : ((forvar330 != forvar330) ~^ $signed(forvar330)))} ?
              reg328[(4'hd):(3'h6)] : reg359[(4'hc):(2'h2)]);
        end
      for (forvar360 = (1'h0); (forvar360 < (1'h0)); forvar360 = (forvar360 + (1'h1)))
        begin
          for (forvar361 = (1'h0); (forvar361 < (1'h1)); forvar361 = (forvar361 + (1'h1)))
            begin
              reg362 <= {(~(&(|reg329[(2'h2):(1'h0)])))};
              reg363 = {(($unsigned(reg310) ^~ {forvar361[(3'h5):(2'h2)]}) << reg310),
                  ((~|($signed((7'h44)) ?
                          (wire295 | (7'h41)) : $unsigned(reg305))) ?
                      reg353[(4'hc):(1'h1)] : reg330[(1'h1):(1'h1)])};
            end
          reg364 <= ((((~|reg312) ? reg305 : (^wire352[(4'ha):(4'h8)])) ?
                  ((~$unsigned(reg329)) ?
                      reg349[(4'h9):(1'h1)] : $signed((wire297 >>> reg353))) : (~|$signed({wire295}))) ?
              {reg333[(4'h9):(2'h3)],
                  (({wire296, reg346} | reg328[(4'h9):(1'h0)]) ?
                      $signed($signed((8'hbf))) : $signed({forvar327}))} : (8'ha6));
        end
    end
  assign wire365 = ($signed(reg306[(3'h6):(3'h6)]) < (~^$unsigned((+wire302[(1'h1):(1'h0)]))));
  assign wire366 = ((reg310[(3'h4):(1'h0)] ~^ ((reg323[(4'hb):(4'h9)] < (8'h9f)) ?
                       (8'hbd) : reg325[(4'h9):(3'h7)])) >= $unsigned((~|$signed((~^reg339)))));
  assign wire367 = $unsigned(((($signed(wire300) ?
                           reg350[(4'h9):(3'h5)] : (forvar345 != reg305)) ?
                       {$signed(forvar347),
                           forvar360[(4'hb):(3'h5)]} : $unsigned(wire342)) > $unsigned($unsigned((^(8'haa))))));
  always
    @(posedge clk) begin
      reg368 <= reg321[(1'h0):(1'h0)];
      reg369 <= forvar327;
    end
  assign wire370 = (+(~|$signed(reg326[(2'h2):(1'h0)])));
  assign wire371 = reg322;
  assign wire372 = (~|reg363);
  assign wire373 = wire298;
  always
    @(posedge clk) begin
      reg374 <= ($unsigned($unsigned((!(^reg305)))) ?
          reg323 : reg330[(1'h1):(1'h0)]);
      if (wire296)
        begin
          reg375 = ($unsigned(wire373) ?
              ($signed((-(reg312 ? reg328 : reg310))) >> reg315) : (8'hb9));
          reg376 <= {($signed("ztI") ?
                  (8'had) : $unsigned((-$signed(reg305))))};
          if (forvar355)
            begin
              reg377 <= $unsigned((wire342[(4'h9):(3'h6)] ?
                  (&(!$unsigned(forvar355))) : ((~$unsigned(reg334)) & (^~(wire352 ?
                      reg368 : wire367)))));
              reg378 = (&("qKL38" ?
                  (($signed(reg333) | "IAwRHm4uHmfhs") >= wire302[(1'h0):(1'h0)]) : reg328[(3'h6):(3'h4)]));
            end
          else
            begin
              reg377 = forvar337[(2'h3):(1'h1)];
              reg378 <= ((~|{reg351[(5'h12):(5'h10)]}) ?
                  reg340[(2'h2):(1'h0)] : $unsigned((((reg335 || wire366) ?
                      $unsigned(wire367) : reg315[(1'h0):(1'h0)]) ^~ $signed((8'hbf)))));
              reg379 <= (((($signed(reg326) ? (8'hbc) : forvar314) ?
                  reg351[(3'h4):(2'h3)] : (~^(^~reg362))) - (~&(((8'hb2) ?
                      reg377 : reg378) ?
                  (-(8'ha3)) : (reg327 ?
                      reg351 : reg344)))) - $unsigned((reg354[(4'hf):(2'h3)] ?
                  $unsigned(reg306) : (reg376 ?
                      ((7'h44) < reg362) : (reg358 ? reg307 : reg330)))));
              reg380 <= (&({"", (8'hb6)} ?
                  (reg325[(2'h3):(1'h0)] ?
                      $signed($unsigned(reg359)) : (((8'ha9) == reg375) ?
                          $unsigned(reg343) : $signed(forvar320))) : $signed((~&reg312))));
              reg381 <= $unsigned($unsigned({reg348}));
            end
          for (forvar382 = (1'h0); (forvar382 < (2'h3)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 <= "UkuLoDMYY";
            end
        end
      else
        begin
          for (forvar375 = (1'h0); (forvar375 < (2'h3)); forvar375 = (forvar375 + (1'h1)))
            begin
              reg376 <= $unsigned((reg310[(2'h3):(2'h3)] <= "cMCPtyZv8XB"));
              reg377 = reg333;
              reg378 = $signed($unsigned(($signed(reg349[(3'h4):(1'h1)]) ?
                  {reg356[(1'h0):(1'h0)]} : ($unsigned(reg306) ?
                      {wire302, forvar355} : reg363[(4'h9):(3'h4)]))));
            end
          reg379 <= $unsigned($signed(reg339[(3'h4):(1'h0)]));
          reg380 <= reg313[(4'h8):(2'h2)];
          if (((("08HMWYbBvzA" || (-reg376)) ?
              $unsigned(forvar347) : {{(forvar360 == (8'haf))},
                  (&forvar382[(3'h5):(1'h1)])}) || wire373[(4'hf):(4'hd)]))
            begin
              reg381 <= {$signed(wire302), (-reg349)};
              reg382 = ((~|(^{wire371})) ?
                  ((!$signed(reg310[(3'h4):(2'h2)])) ?
                      (reg325 ?
                          $unsigned("") : ((|(8'hb9)) ^~ (+reg321))) : forvar309) : {$unsigned((+{reg306}))});
              reg383 <= (forvar318[(2'h3):(2'h3)] ?
                  reg310[(2'h3):(1'h0)] : forvar382[(1'h0):(1'h0)]);
              reg384 <= reg317[(3'h7):(1'h0)];
              reg385 = (~^$unsigned(reg382));
            end
          else
            begin
              reg381 <= ("Vzk3mPs9xH" ?
                  reg334 : $unsigned(($unsigned((&wire302)) ?
                      $unsigned(forvar314) : reg343[(5'h12):(2'h3)])));
              reg382 <= $signed(($signed($unsigned($unsigned(wire301))) ?
                  (("tKyDrMtF5V" ? {(7'h42), reg304} : (^~reg307)) ?
                      $unsigned(forvar375[(2'h2):(1'h0)]) : ({reg313} + reg335[(2'h2):(1'h0)])) : (+{$unsigned(reg375),
                      reg377})));
            end
        end
      reg386 = ($signed((reg327 ?
          reg312 : forvar345[(3'h5):(3'h4)])) ^~ reg364[(2'h2):(2'h2)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module141  (y, clk, wire146, wire145, wire144, wire143, wire142);
  output wire [(32'h5ca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire146;
  input wire [(4'h9):(1'h0)] wire145;
  input wire [(2'h2):(1'h0)] wire144;
  input wire signed [(5'h12):(1'h0)] wire143;
  input wire signed [(4'h8):(1'h0)] wire142;
  reg signed [(3'h4):(1'h0)] reg263 = (1'h0);
  reg [(4'he):(1'h0)] forvar249 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg245 = (1'h0);
  reg [(3'h7):(1'h0)] forvar244 = (1'h0);
  reg [(2'h2):(1'h0)] reg262 = (1'h0);
  reg [(4'h9):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg260 = (1'h0);
  reg [(5'h13):(1'h0)] reg259 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg258 = (1'h0);
  reg [(3'h5):(1'h0)] forvar257 = (1'h0);
  reg [(3'h5):(1'h0)] reg256 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg255 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg254 = (1'h0);
  reg [(5'h12):(1'h0)] reg253 = (1'h0);
  reg signed [(4'he):(1'h0)] reg252 = (1'h0);
  reg [(3'h4):(1'h0)] reg251 = (1'h0);
  reg [(5'h14):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg248 = (1'h0);
  reg [(5'h11):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg246 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar245 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg244 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg243 = (1'h0);
  reg [(4'h9):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg239 = (1'h0);
  reg [(3'h5):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar236 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  reg [(5'h10):(1'h0)] reg234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg233 = (1'h0);
  reg [(5'h15):(1'h0)] reg232 = (1'h0);
  reg [(3'h7):(1'h0)] forvar231 = (1'h0);
  reg [(5'h11):(1'h0)] reg230 = (1'h0);
  reg [(4'h8):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] forvar228 = (1'h0);
  reg [(5'h13):(1'h0)] forvar227 = (1'h0);
  wire [(4'h9):(1'h0)] wire226;
  wire signed [(5'h13):(1'h0)] wire225;
  wire [(5'h15):(1'h0)] wire224;
  wire signed [(2'h2):(1'h0)] wire223;
  wire [(5'h14):(1'h0)] wire222;
  wire signed [(2'h2):(1'h0)] wire221;
  reg signed [(3'h6):(1'h0)] reg220 = (1'h0);
  reg [(5'h15):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg218 = (1'h0);
  reg [(5'h15):(1'h0)] forvar217 = (1'h0);
  reg [(3'h4):(1'h0)] forvar216 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg215 = (1'h0);
  reg [(3'h7):(1'h0)] reg214 = (1'h0);
  reg [(3'h5):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg212 = (1'h0);
  reg [(4'h8):(1'h0)] forvar211 = (1'h0);
  reg [(5'h13):(1'h0)] reg210 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg209 = (1'h0);
  reg [(3'h4):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg206 = (1'h0);
  reg [(4'ha):(1'h0)] reg205 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar204 = (1'h0);
  reg [(5'h13):(1'h0)] reg203 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire202;
  wire [(4'h9):(1'h0)] wire201;
  reg signed [(4'hb):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar195 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg199 = (1'h0);
  reg [(3'h4):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar197 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg196 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg195 = (1'h0);
  reg [(4'ha):(1'h0)] reg194 = (1'h0);
  reg [(5'h15):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg192 = (1'h0);
  reg [(2'h3):(1'h0)] forvar191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg189 = (1'h0);
  reg [(4'ha):(1'h0)] reg188 = (1'h0);
  reg [(4'hc):(1'h0)] reg187 = (1'h0);
  reg [(5'h12):(1'h0)] reg186 = (1'h0);
  reg [(5'h15):(1'h0)] reg185 = (1'h0);
  reg [(3'h5):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg182 = (1'h0);
  reg [(5'h13):(1'h0)] forvar181 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar180 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg179 = (1'h0);
  reg [(4'he):(1'h0)] reg178 = (1'h0);
  reg [(4'hb):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg175 = (1'h0);
  reg [(4'ha):(1'h0)] reg174 = (1'h0);
  reg [(5'h15):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg171 = (1'h0);
  reg [(4'hc):(1'h0)] reg170 = (1'h0);
  reg [(5'h13):(1'h0)] forvar169 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire168;
  reg [(4'h9):(1'h0)] reg167 = (1'h0);
  reg [(5'h15):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg165 = (1'h0);
  reg [(5'h12):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg163 = (1'h0);
  reg [(5'h15):(1'h0)] forvar162 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg161 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg159 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar158 = (1'h0);
  reg [(4'hc):(1'h0)] reg157 = (1'h0);
  reg [(5'h12):(1'h0)] forvar156 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg155 = (1'h0);
  wire [(4'h8):(1'h0)] wire154;
  wire [(2'h3):(1'h0)] wire153;
  wire signed [(3'h4):(1'h0)] wire152;
  wire signed [(4'he):(1'h0)] wire151;
  reg signed [(3'h5):(1'h0)] reg150 = (1'h0);
  reg [(4'hc):(1'h0)] reg149 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire148;
  wire [(4'hc):(1'h0)] wire147;
  assign y = {reg263,
                 forvar249,
                 reg245,
                 forvar244,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 forvar257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 forvar245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 forvar236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 forvar231,
                 reg230,
                 reg229,
                 forvar228,
                 forvar227,
                 wire226,
                 wire225,
                 wire224,
                 wire223,
                 wire222,
                 wire221,
                 reg220,
                 reg219,
                 reg218,
                 forvar217,
                 forvar216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 forvar211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 forvar204,
                 reg203,
                 wire202,
                 wire201,
                 reg200,
                 forvar195,
                 reg199,
                 reg198,
                 forvar197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 forvar181,
                 forvar180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 forvar169,
                 wire168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 forvar162,
                 reg161,
                 reg160,
                 reg159,
                 forvar158,
                 reg157,
                 forvar156,
                 reg155,
                 wire154,
                 wire153,
                 wire152,
                 wire151,
                 reg150,
                 reg149,
                 wire148,
                 wire147,
                 (1'h0)};
  assign wire147 = {$signed(wire145)};
  assign wire148 = $signed((~wire142[(2'h3):(1'h1)]));
  always
    @(posedge clk) begin
      reg149 = (!$signed({(((8'ha8) < wire145) ?
              (~&(8'haa)) : $unsigned(wire142))}));
      reg150 <= ($signed($signed(wire147)) << $unsigned(($unsigned($signed(wire147)) > $unsigned(wire144))));
    end
  assign wire151 = ("gSSQLdKwmh4pshzE" < {$signed(({reg149, wire146} ?
                           wire144 : (|reg149))),
                       $unsigned(wire148)});
  assign wire152 = wire145[(1'h0):(1'h0)];
  assign wire153 = {{(^~wire146), "CQXLd"}};
  assign wire154 = (&((!(+$signed(wire147))) ?
                       $signed((-$unsigned(wire144))) : (^wire144)));
  always
    @(posedge clk) begin
      reg155 <= (wire146 | $unsigned((+(^(wire147 <<< wire146)))));
      for (forvar156 = (1'h0); (forvar156 < (2'h3)); forvar156 = (forvar156 + (1'h1)))
        begin
          reg157 = wire148;
          for (forvar158 = (1'h0); (forvar158 < (3'h4)); forvar158 = (forvar158 + (1'h1)))
            begin
              reg159 = wire147[(3'h7):(2'h2)];
              reg160 <= $unsigned(($signed($unsigned(forvar158)) - (8'hba)));
              reg161 <= wire142;
            end
          for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 = {wire152, (8'hb9)};
              reg164 = reg159;
              reg165 <= (~|(wire154[(2'h2):(1'h0)] || wire152[(2'h2):(1'h1)]));
              reg166 <= wire144;
              reg167 = ({$unsigned({(-(8'ha2))})} != wire154[(3'h4):(2'h3)]);
            end
        end
    end
  assign wire168 = $signed((+((~&forvar156[(1'h1):(1'h1)]) && reg149[(4'hb):(3'h6)])));
  always
    @(posedge clk) begin
      for (forvar169 = (1'h0); (forvar169 < (1'h0)); forvar169 = (forvar169 + (1'h1)))
        begin
          if ({(wire147[(4'hc):(3'h4)] >> (reg149 ?
                  reg149[(3'h6):(1'h1)] : $signed(forvar158)))})
            begin
              reg170 <= $unsigned((8'ha1));
            end
          else
            begin
              reg170 = ($signed(wire146[(4'hd):(2'h3)]) + $signed(({$signed(wire168)} <= wire144)));
              reg171 <= reg163;
              reg172 <= ($unsigned($unsigned("ln2Mm9GUOgkbP")) < reg157[(1'h0):(1'h0)]);
              reg173 = (((8'hb6) && (8'hb9)) ?
                  (!reg167[(4'h8):(3'h4)]) : (reg159 < (~^reg164)));
            end
          reg174 = ({((8'hae) ?
                      $unsigned($unsigned(reg149)) : (wire143 << (~&reg172)))} ?
              $signed($signed($signed(""))) : ((+$unsigned((wire154 ~^ reg155))) ?
                  ((reg155 ? $unsigned(forvar158) : reg171[(3'h7):(3'h5)]) ?
                      ((wire148 >>> wire146) ?
                          (wire148 && (8'ha3)) : reg159[(3'h5):(2'h3)]) : $signed((8'h9d))) : forvar158));
          if ($unsigned((+(wire143[(4'hb):(2'h3)] ?
              ((reg165 ? wire143 : forvar158) ?
                  (!(8'hbf)) : reg164) : reg170))))
            begin
              reg175 <= wire146;
              reg176 <= $signed(reg159[(4'h9):(3'h7)]);
              reg177 <= {reg174};
              reg178 = (^~((reg172 < $signed(reg155)) != $signed(reg160)));
            end
          else
            begin
              reg175 <= $signed($unsigned(((|$unsigned((7'h44))) ?
                  ((reg167 << reg161) > $signed((8'hb4))) : ("ZECR2TeVt4K" ?
                      $signed(wire145) : (|wire144)))));
              reg176 <= (^~((+$signed(reg157[(4'hb):(3'h4)])) || $unsigned($signed(reg157))));
            end
          reg179 <= forvar158[(4'h8):(3'h4)];
        end
      for (forvar180 = (1'h0); (forvar180 < (2'h2)); forvar180 = (forvar180 + (1'h1)))
        begin
          for (forvar181 = (1'h0); (forvar181 < (2'h2)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 <= $unsigned("ASrycCmoIzn0bGAKSDOv");
              reg183 = $signed((reg177 ?
                  (reg166 ?
                      (reg174[(2'h2):(1'h1)] ?
                          $unsigned(reg170) : (reg160 >= reg163)) : $signed((reg173 & forvar162))) : (+(+$unsigned((8'hba))))));
              reg184 = ($signed(($unsigned((&wire146)) <<< (8'ha1))) ?
                  (((forvar162[(4'ha):(3'h6)] == forvar158[(3'h7):(3'h6)]) < (reg173 ?
                      $unsigned(wire146) : $signed(wire168))) && ($signed(reg164) + reg159[(3'h7):(1'h0)])) : $signed((~|((&forvar181) ?
                      (~^(8'ha2)) : wire168))));
            end
          if ((~((wire152[(3'h4):(1'h1)] == (8'ha7)) ~^ reg183)))
            begin
              reg185 <= (&reg166[(4'ha):(1'h1)]);
            end
          else
            begin
              reg185 = ($signed($unsigned((reg177[(4'ha):(3'h4)] ^ $unsigned(reg170)))) ^ {$unsigned(((~^(8'h9d)) ?
                      $signed(reg166) : {reg183}))});
              reg186 <= (($signed(reg157) > reg163[(3'h4):(3'h4)]) ?
                  (8'hac) : (8'h9f));
              reg187 = $unsigned((($signed((8'hb3)) ?
                  $signed(wire143) : $unsigned($signed(wire168))) && $signed($signed((wire154 ^ wire144)))));
              reg188 = reg167;
              reg189 <= $signed($unsigned($unsigned($signed($unsigned((8'hab))))));
            end
        end
      reg190 <= (($signed((^wire142[(1'h0):(1'h0)])) <= ($signed((!reg166)) + $signed($unsigned(wire144)))) ?
          reg160[(1'h1):(1'h1)] : reg176[(5'h15):(4'hc)]);
      for (forvar191 = (1'h0); (forvar191 < (2'h2)); forvar191 = (forvar191 + (1'h1)))
        begin
          reg192 <= (wire151 ?
              ($signed((wire143[(3'h7):(3'h6)] ? reg187 : (^(8'hbc)))) ?
                  $signed((!(reg176 * reg173))) : (reg157[(3'h4):(1'h1)] + $signed(forvar191))) : ((reg163[(4'he):(4'h9)] << $unsigned((&wire147))) ?
                  $signed(reg150[(3'h5):(2'h2)]) : ($signed($signed(forvar180)) ?
                      $unsigned((~^reg171)) : (((8'hbe) ? (8'hab) : reg187) ?
                          (reg157 ?
                              reg189 : (8'hac)) : reg179[(3'h6):(3'h4)]))));
        end
      reg193 <= $unsigned($unsigned($signed(reg179)));
    end
  always
    @(posedge clk) begin
      reg194 <= reg186;
      if ($signed($signed($signed(({(8'h9e), reg188} == $unsigned(reg176))))))
        begin
          reg195 = (^reg183);
          reg196 = reg182[(4'hc):(4'h8)];
          for (forvar197 = (1'h0); (forvar197 < (1'h1)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 <= {(|{(!wire144)})};
            end
          reg199 = $unsigned("tTbRwIsBCb85L");
        end
      else
        begin
          for (forvar195 = (1'h0); (forvar195 < (3'h4)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 = reg199;
            end
          for (forvar197 = (1'h0); (forvar197 < (1'h1)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 <= (reg149 ?
                  (&(reg163 ?
                      ($unsigned((8'hae)) < (|reg188)) : $signed((reg179 ?
                          reg196 : reg193)))) : reg166[(5'h13):(5'h11)]);
              reg199 <= (8'ha7);
              reg200 <= (~|$signed(({(reg189 ?
                      wire168 : wire146)} ~^ $unsigned("fdEr8esxhxlBRsNIBt0"))));
            end
        end
    end
  assign wire201 = reg173[(4'ha):(3'h7)];
  assign wire202 = reg186;
  always
    @(posedge clk) begin
      reg203 <= $signed(reg160);
      for (forvar204 = (1'h0); (forvar204 < (1'h1)); forvar204 = (forvar204 + (1'h1)))
        begin
          if ((($unsigned(((reg172 < reg198) ?
                  wire154[(4'h8):(1'h1)] : $signed(reg203))) ~^ {forvar158,
                  reg173[(4'hf):(2'h3)]}) ?
              ({{(^~forvar162)}} ?
                  "" : reg176[(4'h9):(4'h8)]) : $signed($unsigned((reg192 | reg174)))))
            begin
              reg205 = $unsigned($unsigned({{(reg150 ? (8'hb2) : reg172)}}));
              reg206 <= ($signed(((!$unsigned(wire168)) ?
                      $unsigned((+reg182)) : (^{reg149}))) ?
                  $unsigned($unsigned({reg196})) : reg184);
            end
          else
            begin
              reg205 = (+((8'hbd) ? {reg205} : $unsigned($signed((&reg195)))));
              reg206 = ($unsigned($unsigned(reg200[(4'hb):(3'h7)])) ?
                  "OgcJ1zUYcSp40zvd" : $signed($signed($signed((~(8'hbc))))));
            end
          reg207 <= (((&wire148[(1'h1):(1'h0)]) > (|reg183[(3'h6):(2'h2)])) >= {$unsigned($signed($signed((7'h40)))),
              $unsigned(wire168[(4'hb):(3'h7)])});
          if ((^(!(~|($unsigned(reg183) ?
              (~^(8'hb3)) : reg173[(5'h14):(5'h12)])))))
            begin
              reg208 <= wire148[(1'h0):(1'h0)];
            end
          else
            begin
              reg208 <= reg187[(1'h0):(1'h0)];
              reg209 <= $signed((~&reg165));
            end
          reg210 <= ((~$signed({(reg194 >>> wire144), $unsigned((8'ha4))})) ?
              {reg206,
                  $unsigned($unsigned((reg206 > reg208)))} : (~$signed((((8'ha8) ?
                      forvar156 : wire151) ?
                  $unsigned((7'h43)) : {reg171}))));
          for (forvar211 = (1'h0); (forvar211 < (3'h4)); forvar211 = (forvar211 + (1'h1)))
            begin
              reg212 = (&$signed(((reg157[(4'hc):(1'h0)] || "O3bfP") ?
                  $signed((wire153 == wire148)) : reg171[(4'h8):(3'h5)])));
              reg213 <= $signed(($signed("9K6") * (^~forvar204)));
              reg214 <= reg161;
              reg215 <= reg161[(4'hd):(4'hc)];
            end
        end
      for (forvar216 = (1'h0); (forvar216 < (2'h2)); forvar216 = (forvar216 + (1'h1)))
        begin
          for (forvar217 = (1'h0); (forvar217 < (2'h2)); forvar217 = (forvar217 + (1'h1)))
            begin
              reg218 <= $signed(($unsigned(((~reg193) ~^ {reg161, wire146})) ?
                  {reg161[(4'h8):(3'h6)], reg183} : (~$unsigned(((8'hba) ?
                      reg176 : reg165)))));
              reg219 <= wire153[(1'h0):(1'h0)];
              reg220 <= (reg164[(5'h10):(2'h3)] <= $unsigned(reg149));
            end
        end
    end
  assign wire221 = (^((~&((reg178 || reg213) - $unsigned((8'h9e)))) != reg209[(2'h2):(1'h0)]));
  assign wire222 = wire143;
  assign wire223 = (($signed(reg192) ?
                           {(8'hae),
                               $unsigned((reg208 <= reg173))} : forvar211[(3'h7):(3'h4)]) ?
                       forvar204 : ($unsigned(((reg212 && forvar169) - reg195[(3'h7):(3'h5)])) * ({$signed(wire153),
                               wire142} ?
                           (+(+forvar162)) : {{reg188}})));
  assign wire224 = $signed(wire145);
  assign wire225 = (8'hbd);
  assign wire226 = $signed((~|(wire201 >>> ({reg165,
                       (8'hb3)} + (reg189 < reg159)))));
  always
    @(posedge clk) begin
      for (forvar227 = (1'h0); (forvar227 < (2'h2)); forvar227 = (forvar227 + (1'h1)))
        begin
          for (forvar228 = (1'h0); (forvar228 < (2'h2)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 <= reg195;
              reg230 <= $unsigned(reg205);
            end
          for (forvar231 = (1'h0); (forvar231 < (2'h2)); forvar231 = (forvar231 + (1'h1)))
            begin
              reg232 <= $unsigned({(8'ha9)});
              reg233 = reg200;
              reg234 <= {$unsigned($signed(reg220)),
                  ((-(-reg157[(1'h1):(1'h1)])) | $unsigned((^~forvar169[(3'h6):(1'h0)])))};
              reg235 <= reg174[(1'h0):(1'h0)];
            end
          for (forvar236 = (1'h0); (forvar236 < (2'h3)); forvar236 = (forvar236 + (1'h1)))
            begin
              reg237 = $signed(reg193[(5'h11):(4'ha)]);
              reg238 = $unsigned(reg206[(4'h8):(3'h4)]);
              reg239 <= forvar227;
              reg240 <= reg183[(3'h7):(3'h4)];
              reg241 = $unsigned($unsigned($unsigned(reg179)));
            end
          reg242 <= reg206[(3'h5):(2'h2)];
        end
      reg243 <= (forvar191 ?
          ((($signed((8'ha6)) >= $signed(reg159)) ^~ $signed($unsigned(reg172))) ?
              ($unsigned((wire168 ? reg186 : reg198)) ?
                  (((8'ha5) ? reg176 : wire221) | (reg212 ?
                      reg184 : (8'hbe))) : reg189[(3'h5):(3'h5)]) : (8'ha0)) : reg159);
    end
  always
    @(posedge clk) begin
      if ((~|$signed(wire143)))
        begin
          reg244 = ($signed(reg192) && (^~reg189[(1'h0):(1'h0)]));
          for (forvar245 = (1'h0); (forvar245 < (1'h0)); forvar245 = (forvar245 + (1'h1)))
            begin
              reg246 <= $signed(((reg233 > (8'hba)) << reg210));
            end
          if ($unsigned(reg179[(3'h4):(2'h2)]))
            begin
              reg247 <= $signed($unsigned(reg210));
              reg248 <= reg166[(5'h13):(3'h7)];
              reg249 = reg190[(3'h6):(3'h6)];
              reg250 = $unsigned($signed(($unsigned((forvar245 | reg193)) * $unsigned((reg160 ?
                  reg248 : reg167)))));
            end
          else
            begin
              reg247 = ($signed((((~^reg172) ?
                          (wire225 & wire201) : $unsigned(reg230)) ?
                      reg184 : (|((8'h9d) <= reg157)))) ?
                  reg165[(3'h6):(3'h4)] : $unsigned($unsigned(((wire221 ?
                          reg176 : wire154) ?
                      reg176 : $unsigned(reg157)))));
              reg248 <= (8'hb0);
              reg249 <= reg165;
              reg250 <= reg210[(5'h13):(4'he)];
              reg251 <= {$unsigned($unsigned({wire224}))};
            end
          if ((8'hbc))
            begin
              reg252 <= $signed($signed(($signed((reg187 <<< wire154)) ?
                  $signed(forvar195) : $unsigned(((8'ha4) ?
                      reg242 : reg241)))));
              reg253 <= (~^reg209);
              reg254 = "";
              reg255 <= reg198[(1'h0):(1'h0)];
              reg256 = reg252;
            end
          else
            begin
              reg252 = forvar228[(1'h0):(1'h0)];
              reg253 <= (|((reg233[(4'hd):(4'hd)] ? (8'hb5) : (~^reg206)) ?
                  reg150[(2'h2):(1'h0)] : ({reg230} ?
                      reg207[(4'ha):(3'h5)] : reg244)));
            end
          for (forvar257 = (1'h0); (forvar257 < (2'h2)); forvar257 = (forvar257 + (1'h1)))
            begin
              reg258 <= forvar169[(4'hb):(1'h0)];
              reg259 <= (~|(8'ha0));
              reg260 <= (reg255 ? $unsigned(reg232) : $unsigned((8'ha5)));
              reg261 = $signed($unsigned($unsigned(reg255[(3'h7):(1'h1)])));
              reg262 = (reg175 ? forvar211 : wire226);
            end
        end
      else
        begin
          for (forvar244 = (1'h0); (forvar244 < (2'h3)); forvar244 = (forvar244 + (1'h1)))
            begin
              reg245 <= ($signed($unsigned((-{(8'hbb)}))) != reg237[(3'h7):(3'h6)]);
              reg246 <= (8'h9c);
              reg247 = reg213[(2'h2):(1'h1)];
            end
          if ($unsigned($signed((+(~&"KZK")))))
            begin
              reg248 <= $unsigned((~$signed(forvar211[(2'h2):(1'h0)])));
            end
          else
            begin
              reg248 = $signed(((^({wire225} ?
                  $unsigned(reg241) : reg235[(4'he):(2'h3)])) ^~ forvar245));
            end
          for (forvar249 = (1'h0); (forvar249 < (1'h0)); forvar249 = (forvar249 + (1'h1)))
            begin
              reg250 <= $signed((~^(({reg192} ?
                      reg261 : ((8'hb5) ? (8'haa) : (8'hba))) ?
                  ((wire226 && (8'hb1)) ?
                      $unsigned((8'hbe)) : $signed(reg238)) : (&$signed(reg242)))));
            end
        end
      reg263 <= ($signed(reg195[(2'h3):(1'h1)]) || (+(forvar211 ^ ($signed(wire143) ?
          $signed(reg210) : $signed(forvar216)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module832
#( parameter param925 = {(~&(((~&(8'h9f)) ? (8'ha1) : (~(8'ha7))) > {((8'h9e) >> (8'ha7))})), ((^((&(7'h42)) - ((8'hbe) >>> (7'h42)))) - {{(~(8'ha9))}, ((7'h42) ? (!(8'ha4)) : ((8'h9f) >= (8'hb2)))})} )
(y, clk, wire836, wire835, wire834, wire833);
  output wire [(32'h444):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire836;
  input wire signed [(5'h11):(1'h0)] wire835;
  input wire [(4'h9):(1'h0)] wire834;
  input wire signed [(4'ha):(1'h0)] wire833;
  wire [(5'h12):(1'h0)] wire924;
  reg signed [(3'h5):(1'h0)] reg923 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg922 = (1'h0);
  reg [(4'h9):(1'h0)] reg921 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg920 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg919 = (1'h0);
  reg signed [(4'he):(1'h0)] reg918 = (1'h0);
  reg [(5'h11):(1'h0)] forvar917 = (1'h0);
  reg [(4'he):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg915 = (1'h0);
  reg [(2'h3):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar913 = (1'h0);
  reg signed [(4'he):(1'h0)] reg912 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar911 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg910 = (1'h0);
  reg [(5'h15):(1'h0)] reg909 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg908 = (1'h0);
  reg [(4'hf):(1'h0)] reg907 = (1'h0);
  reg [(5'h13):(1'h0)] reg906 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar905 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire904;
  reg signed [(4'hc):(1'h0)] reg903 = (1'h0);
  reg [(3'h5):(1'h0)] forvar902 = (1'h0);
  reg [(2'h3):(1'h0)] reg901 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar899 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg898 = (1'h0);
  reg [(5'h10):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg895 = (1'h0);
  reg [(4'h9):(1'h0)] reg894 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg892 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg891 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar890 = (1'h0);
  reg [(5'h12):(1'h0)] reg889 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar887 = (1'h0);
  wire [(3'h5):(1'h0)] wire886;
  wire signed [(4'hc):(1'h0)] wire885;
  reg [(5'h10):(1'h0)] reg884 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg883 = (1'h0);
  reg [(5'h15):(1'h0)] reg882 = (1'h0);
  reg [(5'h14):(1'h0)] forvar881 = (1'h0);
  reg [(5'h11):(1'h0)] reg880 = (1'h0);
  reg [(4'hf):(1'h0)] reg879 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg878 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar877 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar876 = (1'h0);
  reg [(4'hc):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg873 = (1'h0);
  reg [(4'ha):(1'h0)] reg872 = (1'h0);
  reg [(5'h12):(1'h0)] reg871 = (1'h0);
  reg [(4'h8):(1'h0)] reg870 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg869 = (1'h0);
  reg [(5'h15):(1'h0)] reg868 = (1'h0);
  reg [(3'h6):(1'h0)] reg867 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar866 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar865 = (1'h0);
  reg [(4'hd):(1'h0)] reg864 = (1'h0);
  reg [(5'h11):(1'h0)] reg863 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar862 = (1'h0);
  reg [(5'h15):(1'h0)] reg861 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg860 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg859 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg858 = (1'h0);
  reg [(2'h3):(1'h0)] reg857 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg856 = (1'h0);
  reg [(4'hb):(1'h0)] forvar855 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg854 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg853 = (1'h0);
  reg [(3'h5):(1'h0)] reg852 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar851 = (1'h0);
  reg [(4'hb):(1'h0)] forvar850 = (1'h0);
  reg [(5'h11):(1'h0)] reg849 = (1'h0);
  wire [(5'h13):(1'h0)] wire848;
  reg signed [(3'h7):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg845 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg844 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg843 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg842 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg841 = (1'h0);
  reg [(3'h7):(1'h0)] reg840 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg839 = (1'h0);
  reg [(5'h13):(1'h0)] reg838 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire837;
  assign y = {wire924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 forvar917,
                 reg916,
                 reg915,
                 reg914,
                 forvar913,
                 reg912,
                 forvar911,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg906,
                 forvar905,
                 wire904,
                 reg903,
                 forvar902,
                 reg901,
                 reg900,
                 forvar899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 forvar893,
                 reg892,
                 reg891,
                 forvar890,
                 reg889,
                 reg888,
                 forvar887,
                 wire886,
                 wire885,
                 reg884,
                 reg883,
                 reg882,
                 forvar881,
                 reg880,
                 reg879,
                 reg878,
                 forvar877,
                 forvar876,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 forvar866,
                 forvar865,
                 reg864,
                 reg863,
                 forvar862,
                 reg861,
                 reg860,
                 reg859,
                 reg858,
                 reg857,
                 reg856,
                 forvar855,
                 reg854,
                 reg853,
                 reg852,
                 forvar851,
                 forvar850,
                 reg849,
                 wire848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg839,
                 reg838,
                 wire837,
                 (1'h0)};
  assign wire837 = wire834;
  always
    @(posedge clk) begin
      reg838 = $signed(($unsigned(wire834) >>> (wire835 ?
          ($signed(wire836) > (8'ha5)) : wire837)));
      if ((((~&$unsigned($unsigned(wire835))) > $unsigned($unsigned(reg838))) > (-"gayC17GN")))
        begin
          if ($unsigned((-wire835[(4'he):(4'hb)])))
            begin
              reg839 = $signed($signed(($unsigned((^~wire836)) || wire833)));
            end
          else
            begin
              reg839 = ($signed((^({wire836, reg838} ?
                  $unsigned(reg838) : $signed(wire836)))) | wire836);
            end
          if (($signed(wire836[(1'h1):(1'h0)]) && (reg839[(2'h2):(1'h1)] != wire833)))
            begin
              reg840 <= (wire837[(3'h5):(3'h5)] << (((wire834[(3'h4):(3'h4)] ^~ $signed(wire834)) <<< (~^(wire833 || reg838))) ~^ wire833[(1'h1):(1'h1)]));
              reg841 <= wire833;
              reg842 = (-(~^$signed($signed("NySBhVoT7QFkKt"))));
              reg843 = (~|(reg838 ^~ reg839));
              reg844 <= (($signed($signed($unsigned(reg841))) << {(wire836 || (^~reg841)),
                      (wire837 != (reg842 ? reg842 : wire835))}) ?
                  reg843[(1'h0):(1'h0)] : $signed({($unsigned(reg840) && "i")}));
            end
          else
            begin
              reg840 <= wire833;
              reg841 <= (($unsigned((^reg842[(1'h0):(1'h0)])) << $signed(reg839)) <<< reg840[(1'h1):(1'h0)]);
              reg842 <= {$signed(wire835[(5'h10):(4'he)]),
                  $signed(("8Zw" > $unsigned($unsigned(wire837))))};
              reg843 <= (wire837[(4'hd):(3'h5)] & "stFnq0TG");
            end
          reg845 = $signed((!($signed((reg844 < reg839)) ?
              (8'hab) : ({wire834, reg838} << {(8'hba)}))));
          reg846 <= $signed(((!wire835) == {$unsigned(reg839[(2'h3):(2'h3)]),
              (((7'h43) && (8'ha6)) ?
                  (reg845 ? reg839 : reg840) : reg838[(4'he):(3'h6)])}));
        end
      else
        begin
          if (reg845)
            begin
              reg839 = $unsigned((~|$unsigned(reg838)));
            end
          else
            begin
              reg839 <= (reg843 ?
                  reg838 : ({wire833,
                      {(+reg842),
                          (reg838 - (8'ha9))}} & (~^wire833[(3'h7):(3'h5)])));
              reg840 = (reg838[(4'hc):(2'h3)] ^~ wire833);
              reg841 = ({$unsigned((~^reg844))} != $signed($signed(reg842)));
            end
          reg842 = ($signed($unsigned(((reg845 >= reg844) ?
              $signed(reg846) : reg845))) * $unsigned((^reg845[(3'h5):(2'h2)])));
        end
      reg847 <= $signed(($unsigned(reg844[(1'h1):(1'h0)]) >> (^(wire835 ?
          reg843 : ((7'h42) + wire835)))));
    end
  assign wire848 = (!{$unsigned(reg843),
                       ((reg846 ? reg846 : reg846) && reg846)});
  always
    @(posedge clk) begin
      reg849 = reg845;
      for (forvar850 = (1'h0); (forvar850 < (1'h0)); forvar850 = (forvar850 + (1'h1)))
        begin
          for (forvar851 = (1'h0); (forvar851 < (2'h2)); forvar851 = (forvar851 + (1'h1)))
            begin
              reg852 <= wire836;
              reg853 <= ($signed($unsigned(reg852[(2'h2):(1'h0)])) ?
                  {$signed((~^reg844[(4'h8):(3'h7)]))} : "A4bdIvRM4B7");
              reg854 = ($unsigned(((((8'hb8) >> wire837) ?
                  (|reg840) : (~reg849)) >>> $signed(reg847[(3'h4):(2'h2)]))) ^~ (^(8'hbf)));
            end
          for (forvar855 = (1'h0); (forvar855 < (1'h0)); forvar855 = (forvar855 + (1'h1)))
            begin
              reg856 <= reg839;
              reg857 = (reg852 ? "JT4iszQoh" : (~{{forvar851}, reg845}));
              reg858 <= (!({(^{forvar855}), $signed($unsigned(forvar855))} ?
                  ($unsigned($signed(reg841)) > $signed((-wire837))) : reg843));
              reg859 <= (-(reg849[(3'h7):(3'h7)] ?
                  ((reg856[(1'h0):(1'h0)] + (reg841 ? reg857 : reg846)) ?
                      $unsigned($signed(forvar850)) : "PMGKdqQKMzB") : $signed(((^reg842) ?
                      wire834 : reg841))));
            end
          reg860 = (^~forvar851);
          reg861 = wire837[(3'h5):(1'h0)];
          for (forvar862 = (1'h0); (forvar862 < (1'h1)); forvar862 = (forvar862 + (1'h1)))
            begin
              reg863 <= $signed(((($signed(reg852) ?
                          (!(8'hb0)) : ((7'h41) && reg852)) ?
                      $signed($signed(reg849)) : $signed($signed(forvar862))) ?
                  wire836 : wire834));
              reg864 = reg840[(1'h1):(1'h0)];
            end
        end
      for (forvar865 = (1'h0); (forvar865 < (3'h4)); forvar865 = (forvar865 + (1'h1)))
        begin
          for (forvar866 = (1'h0); (forvar866 < (3'h4)); forvar866 = (forvar866 + (1'h1)))
            begin
              reg867 = $signed((~|wire834));
              reg868 = $signed(reg845);
              reg869 <= reg845;
              reg870 = (~|reg838);
              reg871 <= reg860[(2'h2):(1'h1)];
            end
          if ((~|reg840[(3'h6):(3'h5)]))
            begin
              reg872 <= (~^reg847[(2'h3):(1'h1)]);
              reg873 = ($signed(reg871[(4'h9):(1'h1)]) ?
                  (-{reg870, reg860}) : {(reg849 ?
                          ("G36JvLfThYd" ?
                              (+reg842) : $signed(reg864)) : $signed((forvar850 == wire834)))});
              reg874 <= (reg854[(3'h6):(2'h3)] ?
                  {$signed((-forvar862[(2'h3):(2'h3)])),
                      (((^~(8'ha8)) ?
                          reg870[(2'h3):(1'h1)] : $signed(reg858)) - forvar865[(3'h7):(2'h3)])} : $unsigned(reg856));
            end
          else
            begin
              reg872 = reg871;
              reg873 <= (reg854 != forvar865[(3'h7):(1'h0)]);
              reg874 = $signed(((8'hb2) ?
                  (+$signed(wire834)) : ({$unsigned(wire833),
                      (|(8'haf))} != $unsigned(reg867[(1'h0):(1'h0)]))));
              reg875 <= $signed(reg872);
            end
        end
      for (forvar876 = (1'h0); (forvar876 < (2'h2)); forvar876 = (forvar876 + (1'h1)))
        begin
          for (forvar877 = (1'h0); (forvar877 < (2'h2)); forvar877 = (forvar877 + (1'h1)))
            begin
              reg878 <= {$signed(wire833[(4'h9):(2'h2)]),
                  $signed({(reg843 ?
                          reg861[(4'ha):(2'h2)] : (forvar851 ?
                              reg853 : (7'h42))),
                      (^(reg841 ? reg856 : reg875))})};
              reg879 = (reg858[(1'h1):(1'h0)] != $unsigned((!(reg859[(2'h2):(2'h2)] ?
                  reg863[(3'h4):(1'h0)] : (reg856 ? reg843 : (8'ha4))))));
            end
          reg880 <= reg857;
          for (forvar881 = (1'h0); (forvar881 < (2'h3)); forvar881 = (forvar881 + (1'h1)))
            begin
              reg882 = "yJxP9zMgn";
            end
          reg883 <= $signed(reg872[(2'h2):(1'h0)]);
          reg884 = {reg880};
        end
    end
  assign wire885 = reg846;
  assign wire886 = reg838;
  always
    @(posedge clk) begin
      for (forvar887 = (1'h0); (forvar887 < (3'h4)); forvar887 = (forvar887 + (1'h1)))
        begin
          reg888 = (+{((reg869 ?
                      (forvar851 ? wire835 : wire835) : (wire837 ?
                          (8'hb6) : reg859)) ?
                  $signed(reg868[(4'h9):(4'h8)]) : reg873[(2'h3):(2'h3)])});
          reg889 = $unsigned($signed(reg873));
          for (forvar890 = (1'h0); (forvar890 < (2'h3)); forvar890 = (forvar890 + (1'h1)))
            begin
              reg891 = (~(~reg859[(1'h0):(1'h0)]));
              reg892 <= $signed(({reg863} << reg852));
            end
          for (forvar893 = (1'h0); (forvar893 < (3'h4)); forvar893 = (forvar893 + (1'h1)))
            begin
              reg894 <= (reg844[(4'h8):(4'h8)] * (~&{$signed((+wire848))}));
              reg895 <= ($signed($signed($unsigned(((8'had) ?
                      reg864 : reg892)))) ?
                  $signed(reg869[(1'h1):(1'h1)]) : reg882[(5'h14):(3'h5)]);
              reg896 = {($signed($unsigned((reg874 ?
                      reg884 : (7'h42)))) != $signed(reg858))};
              reg897 = reg894[(1'h1):(1'h1)];
              reg898 = $unsigned(reg870);
            end
          for (forvar899 = (1'h0); (forvar899 < (2'h3)); forvar899 = (forvar899 + (1'h1)))
            begin
              reg900 = ($signed(forvar862[(1'h1):(1'h1)]) < "0ODyZLnWA");
              reg901 = $signed(($signed(reg869[(2'h2):(1'h1)]) ^~ $unsigned($signed(forvar881[(5'h11):(4'hf)]))));
            end
        end
      for (forvar902 = (1'h0); (forvar902 < (1'h1)); forvar902 = (forvar902 + (1'h1)))
        begin
          reg903 <= $signed((-{reg842[(2'h2):(1'h1)], reg841}));
        end
    end
  assign wire904 = $unsigned(("" & (&forvar887[(2'h3):(1'h1)])));
  always
    @(posedge clk) begin
      for (forvar905 = (1'h0); (forvar905 < (1'h1)); forvar905 = (forvar905 + (1'h1)))
        begin
          if ($unsigned(wire835))
            begin
              reg906 = $signed((~(((reg883 | reg895) ?
                      $unsigned(reg868) : ((8'hb9) ? reg840 : reg900)) ?
                  reg853 : forvar855)));
              reg907 <= $unsigned(reg880);
            end
          else
            begin
              reg906 <= ((&({{reg843}, $signed(reg896)} ?
                      (((8'hbf) - reg898) ?
                          reg852 : (reg856 >> reg898)) : (~&forvar893))) ?
                  (($signed(reg906[(2'h3):(2'h2)]) ?
                          $signed((reg869 ? (8'hb3) : forvar893)) : ({reg853,
                                  reg906} ?
                              (reg897 <<< wire886) : $signed(forvar865))) ?
                      $unsigned((reg860[(3'h5):(1'h0)] ?
                          forvar893 : (~^reg860))) : {{reg880[(3'h6):(3'h5)],
                              reg847[(1'h0):(1'h0)]}}) : reg841[(1'h1):(1'h1)]);
              reg907 <= "hSJ";
              reg908 <= ($signed($signed(reg854)) ?
                  $signed((7'h42)) : $unsigned($signed({(~&forvar850),
                      (reg900 ? reg852 : reg903)})));
            end
          reg909 <= (~&(($unsigned(forvar876) ?
              $unsigned($unsigned(forvar855)) : {$signed(reg908)}) >= $unsigned(reg873[(1'h1):(1'h0)])));
          reg910 = {reg869};
        end
      for (forvar911 = (1'h0); (forvar911 < (1'h0)); forvar911 = (forvar911 + (1'h1)))
        begin
          reg912 <= $unsigned((&$unsigned($unsigned((7'h42)))));
          for (forvar913 = (1'h0); (forvar913 < (2'h2)); forvar913 = (forvar913 + (1'h1)))
            begin
              reg914 = ($unsigned((!reg910)) & (reg879 == reg883));
              reg915 <= ({(((reg889 || (8'ha2)) ?
                          (reg909 ?
                              reg864 : forvar850) : $signed(reg844)) | (~(-forvar865)))} ?
                  (8'ha7) : forvar855);
              reg916 <= reg854;
            end
          for (forvar917 = (1'h0); (forvar917 < (3'h4)); forvar917 = (forvar917 + (1'h1)))
            begin
              reg918 = {(((8'had) || ((~|reg872) ?
                      (^reg869) : (~&reg896))) | {{(reg883 + reg883),
                          (~|(8'hb7))}}),
                  ((!(8'ha2)) ?
                      reg907 : (((forvar887 ?
                          reg871 : reg880) || wire835) || ((8'h9f) != (reg852 <<< reg841))))};
              reg919 = ({$signed(reg906), {(8'hb4), (8'hbc)}} ?
                  $unsigned("RTDgPJHF27Tt") : (reg838[(5'h11):(4'hb)] + (~"CgrM5H")));
              reg920 = reg906[(2'h2):(1'h1)];
              reg921 <= $signed({reg838,
                  ((((8'hba) == (8'hb0)) ?
                      (reg898 ?
                          reg869 : reg889) : $unsigned((8'hb8))) <<< (~&(~|reg920)))});
              reg922 <= reg910[(3'h4):(1'h1)];
            end
        end
      reg923 <= (((reg875 * ((forvar905 >>> reg864) - reg909[(4'hc):(2'h2)])) >= $unsigned({(reg906 ?
              (8'haf) : reg906)})) ^ ((~&wire848) ?
          reg880 : {(((8'hb7) ? reg859 : wire886) <<< ((8'hbf) ?
                  reg897 : wire885)),
              ($signed(forvar865) >>> $signed((8'ha3)))}));
    end
  assign wire924 = reg874;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module645
#( parameter param730 = {({({(8'hb5), (8'hb6)} ? {(8'hab)} : {(8'ha7), (7'h40)}), (8'had)} ? ((((8'hb6) ? (8'ha3) : (8'hb9)) ? (8'ha0) : ((8'hb2) ? (8'hbf) : (8'hb4))) ? ((+(8'ha1)) ? ((8'had) ? (8'h9d) : (7'h44)) : (&(8'hbc))) : (((8'ha6) > (8'hb2)) ? {(8'hb4), (8'h9d)} : ((8'hab) ? (8'hae) : (8'hbd)))) : ({((8'hb2) <<< (8'hb1)), (+(8'h9f))} ? ((^~(7'h44)) <= ((8'hb8) ? (7'h44) : (8'ha4))) : (+((8'hb7) || (8'hbe)))))} )
(y, clk, wire649, wire648, wire647, wire646);
  output wire [(32'h36d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire649;
  input wire [(5'h10):(1'h0)] wire648;
  input wire signed [(4'h8):(1'h0)] wire647;
  input wire signed [(4'h9):(1'h0)] wire646;
  wire signed [(4'hc):(1'h0)] wire729;
  wire signed [(3'h4):(1'h0)] wire728;
  wire [(3'h4):(1'h0)] wire727;
  wire signed [(4'h9):(1'h0)] wire726;
  reg [(2'h2):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg724 = (1'h0);
  reg [(4'hc):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg721 = (1'h0);
  reg [(4'hc):(1'h0)] reg720 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg719 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg717 = (1'h0);
  reg [(4'hd):(1'h0)] reg716 = (1'h0);
  reg [(4'hd):(1'h0)] reg715 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire714;
  wire signed [(5'h15):(1'h0)] wire713;
  wire signed [(3'h4):(1'h0)] wire712;
  wire [(3'h6):(1'h0)] wire711;
  wire [(2'h2):(1'h0)] wire710;
  wire signed [(3'h6):(1'h0)] wire709;
  wire [(4'h8):(1'h0)] wire708;
  reg [(4'h8):(1'h0)] reg707 = (1'h0);
  wire [(5'h12):(1'h0)] wire706;
  wire signed [(4'hf):(1'h0)] wire705;
  reg signed [(3'h5):(1'h0)] reg704 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire703;
  reg [(3'h4):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg701 = (1'h0);
  reg [(4'hc):(1'h0)] reg700 = (1'h0);
  reg [(2'h2):(1'h0)] reg699 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg698 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg697 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg695 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg694 = (1'h0);
  reg [(5'h10):(1'h0)] reg693 = (1'h0);
  reg [(4'hd):(1'h0)] reg692 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar691 = (1'h0);
  reg [(4'hf):(1'h0)] reg690 = (1'h0);
  reg [(4'h8):(1'h0)] forvar689 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg688 = (1'h0);
  reg [(5'h11):(1'h0)] reg687 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg685 = (1'h0);
  reg [(4'he):(1'h0)] reg684 = (1'h0);
  reg [(2'h2):(1'h0)] reg683 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg681 = (1'h0);
  reg [(3'h4):(1'h0)] reg680 = (1'h0);
  reg [(2'h2):(1'h0)] reg679 = (1'h0);
  reg [(4'h8):(1'h0)] reg678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg677 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar675 = (1'h0);
  reg [(4'h9):(1'h0)] forvar659 = (1'h0);
  reg [(4'h9):(1'h0)] reg655 = (1'h0);
  reg [(3'h7):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg672 = (1'h0);
  reg [(2'h2):(1'h0)] reg671 = (1'h0);
  reg [(4'h9):(1'h0)] reg670 = (1'h0);
  reg [(5'h15):(1'h0)] reg669 = (1'h0);
  reg [(5'h13):(1'h0)] forvar668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg667 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar666 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg664 = (1'h0);
  reg [(3'h7):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg662 = (1'h0);
  reg [(4'ha):(1'h0)] reg661 = (1'h0);
  reg [(5'h14):(1'h0)] reg660 = (1'h0);
  reg [(3'h5):(1'h0)] reg659 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg658 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg657 = (1'h0);
  reg [(5'h10):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar655 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg654 = (1'h0);
  reg [(5'h14):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg652 = (1'h0);
  reg [(4'h8):(1'h0)] forvar651 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar650 = (1'h0);
  assign y = {wire729,
                 wire728,
                 wire727,
                 wire726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 wire714,
                 wire713,
                 wire712,
                 wire711,
                 wire710,
                 wire709,
                 wire708,
                 reg707,
                 wire706,
                 wire705,
                 reg704,
                 wire703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 forvar691,
                 reg690,
                 forvar689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 forvar682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 forvar675,
                 forvar659,
                 reg655,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 forvar668,
                 reg667,
                 forvar666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 reg658,
                 reg657,
                 reg656,
                 forvar655,
                 reg654,
                 reg653,
                 reg652,
                 forvar651,
                 forvar650,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar650 = (1'h0); (forvar650 < (3'h4)); forvar650 = (forvar650 + (1'h1)))
        begin
          for (forvar651 = (1'h0); (forvar651 < (2'h3)); forvar651 = (forvar651 + (1'h1)))
            begin
              reg652 <= {$unsigned((+(forvar651 ?
                      wire646 : (forvar651 >= wire649))))};
            end
          if (wire649[(4'hf):(3'h6)])
            begin
              reg653 <= (~&($signed((^~{reg652})) && {{(reg652 ?
                          wire649 : forvar650),
                      (forvar651 >>> wire649)},
                  ("2g2RznnXX4GDZHUrD" ? wire647 : (-forvar651))}));
              reg654 <= {forvar651,
                  ($unsigned((forvar650[(4'h8):(4'h8)] == (|reg652))) ?
                      ((7'h43) ?
                          wire646[(3'h4):(2'h2)] : $signed("itk")) : reg652[(1'h1):(1'h1)])};
            end
          else
            begin
              reg653 = reg653[(4'ha):(4'h9)];
            end
        end
      if ({reg654[(3'h6):(3'h6)], reg654[(3'h7):(3'h4)]})
        begin
          for (forvar655 = (1'h0); (forvar655 < (1'h1)); forvar655 = (forvar655 + (1'h1)))
            begin
              reg656 <= (8'ha1);
              reg657 <= {(+({(^~forvar655)} + $unsigned((~reg656))))};
              reg658 <= (($unsigned((^$unsigned(reg657))) ?
                      ($unsigned(wire649) >> ($unsigned(reg652) + (&wire647))) : (((reg656 ?
                                  wire649 : (8'hb7)) ?
                              {wire648} : reg652[(1'h0):(1'h0)]) ?
                          (reg653 ?
                              (wire646 ?
                                  forvar655 : wire647) : $unsigned(forvar655)) : (~|(~wire647)))) ?
                  ({(~^(^~wire647))} != $signed(wire649)) : {(($signed(forvar650) >= $signed(forvar651)) ?
                          $unsigned((reg652 ?
                              wire649 : wire646)) : $unsigned((forvar650 != forvar651))),
                      ((forvar655[(4'hd):(2'h3)] ^~ forvar650[(4'hb):(2'h2)]) ?
                          ((-reg652) ?
                              {wire646,
                                  reg652} : $signed((8'ha7))) : $signed(reg657))});
              reg659 <= (wire648[(4'hf):(4'hd)] ?
                  ($unsigned((~|(!(8'ha9)))) ?
                      $signed($signed("q0ZbLEyhlziR")) : $unsigned(forvar655[(3'h6):(3'h4)])) : (^$signed(forvar655[(5'h11):(1'h1)])));
              reg660 <= ($signed($signed((^~(+wire648)))) ?
                  reg657 : reg658[(2'h2):(1'h1)]);
            end
          if ($unsigned(reg657[(4'hf):(1'h1)]))
            begin
              reg661 <= $unsigned((~&$unsigned(($unsigned(reg652) ?
                  reg656 : $unsigned(forvar651)))));
              reg662 <= ($unsigned($signed($signed((&wire649)))) ^ forvar651);
              reg663 <= (~|$signed($unsigned(($unsigned(forvar655) != {reg659}))));
              reg664 <= {reg660[(3'h7):(2'h2)],
                  $unsigned(reg658[(2'h2):(1'h0)])};
              reg665 <= (forvar651 ?
                  reg662[(3'h4):(1'h0)] : ($unsigned(((+reg659) ?
                      $signed(forvar651) : {reg663})) - $unsigned($unsigned((reg664 ^ forvar650)))));
            end
          else
            begin
              reg661 <= $signed((~|$signed(forvar650[(4'ha):(3'h5)])));
              reg662 = ($unsigned((&$unsigned({reg662}))) || $unsigned({($unsigned((8'hb6)) ?
                      reg652[(2'h2):(1'h1)] : reg657[(4'h9):(3'h5)])}));
              reg663 = ((~(8'hb6)) << reg659[(1'h1):(1'h1)]);
            end
          for (forvar666 = (1'h0); (forvar666 < (2'h3)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 = ($signed(wire647) ?
                  forvar666[(3'h6):(1'h1)] : (+forvar655));
            end
          for (forvar668 = (1'h0); (forvar668 < (3'h4)); forvar668 = (forvar668 + (1'h1)))
            begin
              reg669 <= (-reg654);
              reg670 = $unsigned(({(^((8'ha6) ?
                      wire647 : forvar666))} <<< (forvar651 > ((forvar668 ?
                  forvar655 : forvar651) <= (reg661 ? reg667 : reg665)))));
              reg671 <= $unsigned(reg663);
            end
          if (($unsigned($signed("vqJCE6")) ? (+reg654) : (~^"WK24")))
            begin
              reg672 = {"0brtW", reg669[(4'hd):(4'hc)]};
              reg673 <= (($unsigned({(8'hb1)}) ?
                      reg669 : $signed((^{(8'hba), reg669}))) ?
                  reg656 : (((reg660 & (8'ha8)) ~^ (+(-forvar668))) * reg661[(1'h0):(1'h0)]));
            end
          else
            begin
              reg672 <= forvar650[(1'h1):(1'h1)];
              reg673 = (reg654 ? $signed((8'ha7)) : reg661[(1'h0):(1'h0)]);
              reg674 <= reg660;
            end
        end
      else
        begin
          reg655 <= (reg656[(5'h10):(5'h10)] ^ $signed($unsigned((+{(8'haa)}))));
          reg656 <= $signed("ewKE1NMboutTW5aXi5JX");
          reg657 = (reg657 ?
              {$signed(forvar655),
                  forvar655[(5'h10):(4'hf)]} : ((~^((reg672 ^~ forvar666) ?
                  (|reg661) : reg667[(1'h1):(1'h1)])) * (reg658[(2'h2):(1'h1)] * ((reg672 ?
                      reg661 : reg658) ?
                  reg673 : reg655[(1'h0):(1'h0)]))));
          reg658 <= (reg667 < (~$signed($signed(reg657))));
          for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = ($signed(reg654) != $unsigned({(~(reg661 ?
                      reg652 : reg652)),
                  (wire649 ?
                      ((8'hab) ?
                          forvar655 : forvar666) : reg664[(1'h0):(1'h0)])}));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar675 = (1'h0); (forvar675 < (2'h3)); forvar675 = (forvar675 + (1'h1)))
        begin
          reg676 = ((+reg653[(3'h5):(3'h4)]) + (reg658[(1'h1):(1'h0)] | wire648));
          if (((~^$signed(forvar668[(2'h2):(2'h2)])) ?
              $signed(((((8'ha8) ? reg672 : reg669) >= (reg654 ?
                      reg655 : reg655)) ?
                  (!(reg670 ?
                      reg657 : reg673)) : {(|reg674)})) : $signed((~^($signed(forvar651) ?
                  $signed(reg670) : (~reg664))))))
            begin
              reg677 = $signed($signed((+$signed($signed(wire646)))));
              reg678 = $signed((({$unsigned(reg664), (&forvar668)} ?
                      ((reg655 ?
                          reg657 : reg657) - $unsigned(wire648)) : $unsigned((reg674 ^~ reg653))) ?
                  ((8'h9d) ?
                      $unsigned(forvar650[(4'hf):(1'h0)]) : ({(7'h41),
                          reg656} << $unsigned(reg664))) : ($signed($unsigned(reg672)) ?
                      (&(~^reg665)) : $signed(reg669))));
            end
          else
            begin
              reg677 = forvar668;
              reg678 <= $unsigned(forvar651);
              reg679 <= (((($unsigned((8'hbf)) > (reg676 > wire646)) ?
                      ($signed(wire647) & $signed(wire647)) : (7'h43)) ?
                  (forvar655 ?
                      $signed((forvar666 ?
                          reg674 : reg652)) : $unsigned("Vt10CisoSRXQsDN")) : (~{(reg678 << reg656)})) & (~^(-{(forvar650 || reg665),
                  $signed(reg662)})));
              reg680 <= reg678[(2'h3):(2'h3)];
              reg681 <= reg659;
            end
          for (forvar682 = (1'h0); (forvar682 < (3'h4)); forvar682 = (forvar682 + (1'h1)))
            begin
              reg683 = $unsigned(($signed($unsigned({reg659})) ?
                  (~&$signed((reg655 | reg663))) : reg678));
              reg684 <= {$unsigned(({((7'h42) && reg660)} >> (|(reg663 | reg661)))),
                  reg672[(5'h10):(4'hc)]};
              reg685 <= ($unsigned(($unsigned(reg671[(1'h0):(1'h0)]) ?
                      $signed("QRFBAsMTCQERzn7rH1u") : forvar650)) ?
                  forvar666 : reg653[(4'hf):(3'h4)]);
              reg686 <= ((!reg673[(3'h7):(1'h1)]) ?
                  (7'h44) : (($unsigned(reg683[(2'h2):(1'h0)]) >= $signed(wire649)) ?
                      (~^reg684[(3'h5):(1'h1)]) : (reg684 ?
                          {"Dm", (reg663 && reg659)} : reg681[(4'ha):(3'h5)])));
            end
        end
      reg687 <= reg659[(2'h3):(1'h1)];
      reg688 = reg662;
      for (forvar689 = (1'h0); (forvar689 < (1'h1)); forvar689 = (forvar689 + (1'h1)))
        begin
          reg690 <= $signed(reg653);
          for (forvar691 = (1'h0); (forvar691 < (2'h3)); forvar691 = (forvar691 + (1'h1)))
            begin
              reg692 <= ($signed($unsigned(reg685[(1'h0):(1'h0)])) - ($unsigned(({reg670,
                          reg688} ?
                      (reg681 ? reg658 : reg667) : reg672)) ?
                  ((^(&reg659)) ?
                      ((^forvar659) >>> reg674) : {(reg664 ?
                              wire648 : reg664)}) : (reg672 <<< wire647)));
              reg693 <= $signed((forvar668 && reg658));
              reg694 = reg663[(2'h2):(1'h1)];
              reg695 = reg677;
              reg696 = $unsigned((reg652 ?
                  (wire646 ?
                      reg677 : $signed((-reg657))) : (reg657 || (~(~^forvar650)))));
            end
          reg697 = (reg687[(5'h10):(2'h2)] <= $unsigned(wire649[(4'h8):(1'h1)]));
          if ((forvar675 ?
              (({(-forvar650),
                      forvar659[(2'h2):(1'h0)]} ~^ $unsigned((forvar651 * (8'hb0)))) ?
                  (((reg664 <= reg673) ? (~reg658) : $unsigned(reg679)) ?
                      (+(reg667 + reg671)) : (^~(8'had))) : ($signed((reg696 ^ forvar659)) ?
                      (~|$unsigned(reg693)) : $unsigned((reg661 ?
                          reg656 : reg659)))) : (((+$unsigned((8'hb6))) ^ (~^(|reg658))) ?
                  $signed($signed($unsigned(reg681))) : forvar691)))
            begin
              reg698 = (($signed((((8'hbb) ? (8'hb3) : reg655) ?
                      (reg654 != forvar689) : (reg652 >= reg696))) << ((+(reg659 ?
                          reg669 : wire649)) ?
                      forvar691 : ($signed(reg660) ?
                          (reg688 ? (8'haa) : reg665) : reg693))) ?
                  (($signed(forvar675) && ((&reg656) ~^ (reg693 >>> forvar689))) ?
                      reg690 : {$unsigned($unsigned(reg695)),
                          ((forvar682 ?
                              reg690 : (8'hb5)) >>> $unsigned((8'h9f)))}) : $signed((^forvar691)));
              reg699 <= (wire647 ~^ (~|reg695));
            end
          else
            begin
              reg698 <= (reg686 ?
                  (reg677[(4'h8):(2'h3)] < $signed(reg674)) : $signed(reg679));
              reg699 = ($signed(({(~^forvar659)} || $unsigned((|(8'hb9))))) ?
                  (reg671 ?
                      (+$unsigned((~^reg685))) : reg661) : $signed($signed(($signed(reg679) ?
                      (forvar689 >>> reg687) : $unsigned((7'h44))))));
              reg700 <= ($signed($unsigned(reg663[(3'h7):(3'h4)])) <= reg695);
              reg701 = ($signed(reg664[(1'h0):(1'h0)]) << reg688);
            end
          reg702 <= $signed($signed($unsigned($signed(reg694))));
        end
    end
  assign wire703 = {reg696};
  always
    @(posedge clk) begin
      reg704 = $signed((reg657[(4'hb):(4'hb)] ?
          $unsigned(((reg699 < reg692) ~^ forvar651)) : (~&reg693)));
    end
  assign wire705 = (8'hb6);
  assign wire706 = {$signed(($unsigned(reg667) ?
                           $signed((reg677 ?
                               reg669 : reg653)) : {reg697[(4'h9):(3'h4)],
                               (reg685 - reg696)})),
                       reg660};
  always
    @(posedge clk) begin
      reg707 = $signed(reg656);
    end
  assign wire708 = (reg695 ? (!$unsigned("JkvwNGry")) : reg686);
  assign wire709 = (reg670[(1'h1):(1'h1)] ? reg677[(3'h4):(2'h3)] : forvar689);
  assign wire710 = reg664;
  assign wire711 = {$signed($unsigned((forvar650[(4'hb):(4'h9)] ?
                           (reg667 ^~ reg670) : ((8'hbf) ?
                               forvar666 : reg659))))};
  assign wire712 = reg701[(2'h2):(2'h2)];
  assign wire713 = reg669;
  assign wire714 = ((&reg662[(2'h2):(1'h1)]) ?
                       $signed($unsigned(reg694)) : ($signed(wire708[(4'h8):(2'h2)]) ?
                           $signed(reg698[(1'h1):(1'h0)]) : $signed((((8'ha0) || reg670) ?
                               forvar668[(4'h9):(2'h2)] : {wire711,
                                   wire713}))));
  always
    @(posedge clk) begin
      reg715 <= reg669;
      if ($signed(({((8'hba) ? reg653 : {reg674, wire647}), (8'hbb)} ?
          $unsigned((reg677[(3'h7):(3'h4)] ?
              wire710[(1'h1):(1'h0)] : reg678[(3'h5):(3'h5)])) : {((^~reg653) << (reg676 ^ reg692)),
              reg701})))
        begin
          reg716 <= reg690;
        end
      else
        begin
          reg716 = (~^({$signed(reg655[(4'h8):(1'h1)])} & (~($signed(wire710) ^~ ((8'hb0) ?
              forvar691 : reg690)))));
          reg717 <= (($signed((reg665[(5'h11):(1'h0)] ?
              ((8'ha1) ^~ forvar651) : reg659[(1'h1):(1'h1)])) >> (((reg654 ?
                  wire709 : wire705) ~^ reg681[(2'h3):(1'h1)]) ?
              wire708[(2'h2):(1'h1)] : (reg670 ^~ reg664))) | $signed((-($unsigned(reg658) != $signed((8'hbb))))));
          if (reg654)
            begin
              reg718 <= reg698;
              reg719 = $unsigned(("Bnr" ?
                  (^wire649[(4'h8):(3'h4)]) : $signed(reg652[(1'h1):(1'h0)])));
              reg720 = wire709;
              reg721 <= (|$signed(reg697[(2'h3):(2'h3)]));
            end
          else
            begin
              reg718 = {($unsigned(forvar668[(5'h13):(4'hc)]) < wire708[(3'h6):(2'h3)])};
              reg719 <= (!reg688[(1'h1):(1'h1)]);
              reg720 = reg661[(4'ha):(1'h0)];
            end
          if ($unsigned(wire714))
            begin
              reg722 <= reg694[(2'h3):(1'h0)];
              reg723 <= $unsigned(((~&reg688[(1'h0):(1'h0)]) >> reg680[(1'h1):(1'h1)]));
              reg724 = reg670[(2'h2):(1'h1)];
            end
          else
            begin
              reg722 <= $signed(wire709[(1'h1):(1'h1)]);
              reg723 <= reg721[(3'h4):(2'h3)];
              reg724 = forvar666[(2'h3):(1'h0)];
              reg725 <= $signed((~|reg655[(4'h9):(4'h8)]));
            end
        end
    end
  assign wire726 = $unsigned(((8'hbc) <<< reg699[(2'h2):(1'h0)]));
  assign wire727 = reg683;
  assign wire728 = (reg722[(4'ha):(3'h5)] << $signed(reg721));
  assign wire729 = ({((~{reg716}) > $signed(reg690))} == reg670[(3'h5):(3'h4)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module442
#( parameter param642 = (!((~^(~|(-(8'hac)))) - ({{(8'hb9), (8'ha4)}} + {((7'h44) >> (7'h42))}))) )
(y, clk, wire446, wire445, wire444, wire443);
  output wire [(32'h8b5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire446;
  input wire signed [(3'h5):(1'h0)] wire445;
  input wire signed [(5'h15):(1'h0)] wire444;
  input wire [(4'ha):(1'h0)] wire443;
  wire [(3'h5):(1'h0)] wire641;
  reg [(5'h15):(1'h0)] reg640 = (1'h0);
  reg [(2'h3):(1'h0)] reg639 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg638 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg637 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar636 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg635 = (1'h0);
  reg [(5'h12):(1'h0)] reg634 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg633 = (1'h0);
  reg [(4'hd):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar631 = (1'h0);
  reg [(4'hc):(1'h0)] reg630 = (1'h0);
  reg [(4'hf):(1'h0)] reg629 = (1'h0);
  reg [(3'h5):(1'h0)] reg628 = (1'h0);
  reg [(2'h3):(1'h0)] forvar627 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg626 = (1'h0);
  reg [(4'ha):(1'h0)] reg625 = (1'h0);
  reg [(3'h7):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg623 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar621 = (1'h0);
  reg [(4'he):(1'h0)] reg620 = (1'h0);
  reg [(3'h6):(1'h0)] reg619 = (1'h0);
  reg [(4'he):(1'h0)] forvar618 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg617 = (1'h0);
  reg [(5'h12):(1'h0)] reg616 = (1'h0);
  reg [(4'ha):(1'h0)] reg615 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg613 = (1'h0);
  reg [(4'hc):(1'h0)] forvar612 = (1'h0);
  reg [(3'h4):(1'h0)] reg611 = (1'h0);
  reg [(2'h2):(1'h0)] reg610 = (1'h0);
  reg [(5'h11):(1'h0)] reg609 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg608 = (1'h0);
  reg [(3'h4):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg606 = (1'h0);
  reg [(5'h11):(1'h0)] reg605 = (1'h0);
  reg [(5'h14):(1'h0)] forvar604 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg603 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg598 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg596 = (1'h0);
  reg [(4'ha):(1'h0)] reg602 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg601 = (1'h0);
  reg [(5'h10):(1'h0)] reg600 = (1'h0);
  reg [(4'ha):(1'h0)] reg599 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar598 = (1'h0);
  reg [(3'h4):(1'h0)] reg597 = (1'h0);
  reg [(2'h2):(1'h0)] forvar596 = (1'h0);
  wire [(2'h2):(1'h0)] wire595;
  reg [(5'h12):(1'h0)] forvar589 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg588 = (1'h0);
  reg [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(4'hb):(1'h0)] forvar593 = (1'h0);
  reg [(2'h2):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg591 = (1'h0);
  reg [(3'h6):(1'h0)] reg590 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg589 = (1'h0);
  reg [(4'hf):(1'h0)] forvar588 = (1'h0);
  reg [(3'h7):(1'h0)] reg587 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg586 = (1'h0);
  reg [(5'h14):(1'h0)] reg585 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg584 = (1'h0);
  reg [(4'ha):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar582 = (1'h0);
  reg [(4'h8):(1'h0)] reg581 = (1'h0);
  reg [(4'ha):(1'h0)] reg580 = (1'h0);
  reg [(2'h3):(1'h0)] forvar579 = (1'h0);
  reg [(4'hb):(1'h0)] reg578 = (1'h0);
  reg [(5'h11):(1'h0)] reg577 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg576 = (1'h0);
  reg [(4'h9):(1'h0)] forvar575 = (1'h0);
  reg [(5'h14):(1'h0)] reg574 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg573 = (1'h0);
  reg [(4'hf):(1'h0)] reg572 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar571 = (1'h0);
  reg [(4'hb):(1'h0)] reg570 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg569 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar568 = (1'h0);
  reg [(4'ha):(1'h0)] reg567 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg566 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire565;
  reg [(5'h11):(1'h0)] reg564 = (1'h0);
  reg [(4'hf):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg562 = (1'h0);
  reg [(3'h7):(1'h0)] reg561 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar560 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg559 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg558 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar557 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar556 = (1'h0);
  reg [(4'ha):(1'h0)] forvar554 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar551 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg553 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar552 = (1'h0);
  reg [(3'h6):(1'h0)] reg551 = (1'h0);
  reg [(4'he):(1'h0)] reg550 = (1'h0);
  reg [(5'h10):(1'h0)] forvar549 = (1'h0);
  wire [(5'h15):(1'h0)] wire548;
  reg [(5'h11):(1'h0)] forvar542 = (1'h0);
  reg [(4'h9):(1'h0)] reg540 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar536 = (1'h0);
  reg [(3'h7):(1'h0)] reg547 = (1'h0);
  reg [(2'h2):(1'h0)] forvar546 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg545 = (1'h0);
  reg [(4'h9):(1'h0)] reg544 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg542 = (1'h0);
  reg [(2'h3):(1'h0)] reg541 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar540 = (1'h0);
  reg [(3'h5):(1'h0)] reg539 = (1'h0);
  reg [(4'hd):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg537 = (1'h0);
  reg [(5'h14):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg534 = (1'h0);
  reg [(4'hf):(1'h0)] forvar533 = (1'h0);
  reg [(5'h15):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg530 = (1'h0);
  reg [(5'h14):(1'h0)] reg529 = (1'h0);
  reg [(2'h2):(1'h0)] forvar528 = (1'h0);
  reg [(4'hc):(1'h0)] reg527 = (1'h0);
  reg [(5'h15):(1'h0)] reg526 = (1'h0);
  reg [(3'h4):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg524 = (1'h0);
  reg [(5'h14):(1'h0)] reg523 = (1'h0);
  reg [(3'h5):(1'h0)] forvar522 = (1'h0);
  reg [(5'h14):(1'h0)] reg521 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar519 = (1'h0);
  reg [(4'ha):(1'h0)] reg518 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg517 = (1'h0);
  reg [(4'hb):(1'h0)] reg516 = (1'h0);
  reg [(4'h8):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar514 = (1'h0);
  reg [(4'he):(1'h0)] reg513 = (1'h0);
  reg [(5'h15):(1'h0)] reg512 = (1'h0);
  reg [(3'h5):(1'h0)] reg511 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg510 = (1'h0);
  reg [(5'h10):(1'h0)] reg509 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg508 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar507 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg506 = (1'h0);
  reg [(3'h7):(1'h0)] forvar505 = (1'h0);
  reg [(5'h15):(1'h0)] reg504 = (1'h0);
  wire [(5'h14):(1'h0)] wire503;
  reg [(5'h10):(1'h0)] reg502 = (1'h0);
  reg [(3'h7):(1'h0)] reg501 = (1'h0);
  reg [(3'h4):(1'h0)] reg500 = (1'h0);
  reg [(5'h15):(1'h0)] reg499 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg497 = (1'h0);
  reg [(4'h8):(1'h0)] forvar496 = (1'h0);
  reg [(3'h7):(1'h0)] reg495 = (1'h0);
  reg [(2'h3):(1'h0)] reg494 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar493 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar492 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire491;
  wire signed [(4'hd):(1'h0)] wire490;
  reg signed [(4'h9):(1'h0)] reg489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg [(4'h8):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg486 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg485 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg484 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg483 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar481 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg480 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar479 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg478 = (1'h0);
  reg [(4'hc):(1'h0)] reg477 = (1'h0);
  reg [(3'h5):(1'h0)] reg476 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg475 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar474 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg471 = (1'h0);
  reg [(4'hf):(1'h0)] reg470 = (1'h0);
  reg [(5'h12):(1'h0)] forvar469 = (1'h0);
  reg [(5'h11):(1'h0)] forvar468 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg467 = (1'h0);
  reg [(3'h7):(1'h0)] forvar466 = (1'h0);
  reg [(5'h15):(1'h0)] reg465 = (1'h0);
  reg [(4'h8):(1'h0)] forvar464 = (1'h0);
  reg [(3'h6):(1'h0)] reg463 = (1'h0);
  reg signed [(4'he):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg461 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg460 = (1'h0);
  reg [(3'h7):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg457 = (1'h0);
  reg [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  reg [(4'hb):(1'h0)] reg454 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg453 = (1'h0);
  reg [(5'h10):(1'h0)] forvar452 = (1'h0);
  reg [(2'h2):(1'h0)] forvar451 = (1'h0);
  reg [(4'h9):(1'h0)] reg450 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar449 = (1'h0);
  reg [(4'hf):(1'h0)] forvar448 = (1'h0);
  wire [(4'he):(1'h0)] wire447;
  assign y = {wire641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 forvar636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 forvar631,
                 reg630,
                 reg629,
                 reg628,
                 forvar627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 forvar621,
                 reg620,
                 reg619,
                 forvar618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 forvar612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 forvar604,
                 reg603,
                 reg598,
                 reg596,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 forvar598,
                 reg597,
                 forvar596,
                 wire595,
                 forvar589,
                 reg588,
                 reg594,
                 forvar593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 forvar588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 forvar582,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg577,
                 reg576,
                 forvar575,
                 reg574,
                 reg573,
                 reg572,
                 forvar571,
                 reg570,
                 reg569,
                 forvar568,
                 reg567,
                 reg566,
                 wire565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 forvar560,
                 reg559,
                 reg558,
                 forvar557,
                 forvar556,
                 forvar554,
                 reg552,
                 forvar551,
                 reg555,
                 reg554,
                 reg553,
                 forvar552,
                 reg551,
                 reg550,
                 forvar549,
                 wire548,
                 forvar542,
                 reg540,
                 forvar536,
                 reg547,
                 forvar546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 forvar540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 forvar533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 forvar528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 forvar522,
                 reg521,
                 reg520,
                 forvar519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 forvar507,
                 reg506,
                 forvar505,
                 reg504,
                 wire503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 forvar496,
                 reg495,
                 reg494,
                 forvar493,
                 forvar492,
                 wire491,
                 wire490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 forvar481,
                 reg480,
                 forvar479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 forvar474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 forvar469,
                 forvar468,
                 reg467,
                 forvar466,
                 reg465,
                 forvar464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 forvar452,
                 forvar451,
                 reg450,
                 forvar449,
                 forvar448,
                 wire447,
                 (1'h0)};
  assign wire447 = (~wire444[(3'h6):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar448 = (1'h0); (forvar448 < (2'h3)); forvar448 = (forvar448 + (1'h1)))
        begin
          for (forvar449 = (1'h0); (forvar449 < (2'h2)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 <= ((~&$unsigned(((wire444 ? forvar449 : wire444) ?
                      ((8'hb1) | forvar448) : $signed(forvar448)))) ?
                  $signed($unsigned($signed(wire445))) : (forvar448 >>> {wire443[(1'h0):(1'h0)]}));
            end
        end
      for (forvar451 = (1'h0); (forvar451 < (3'h4)); forvar451 = (forvar451 + (1'h1)))
        begin
          for (forvar452 = (1'h0); (forvar452 < (2'h3)); forvar452 = (forvar452 + (1'h1)))
            begin
              reg453 <= (!(~^$signed($unsigned(forvar448))));
              reg454 <= wire445[(3'h5):(2'h3)];
              reg455 <= (~(wire445[(1'h1):(1'h1)] >>> {((wire446 != reg453) ?
                      wire447 : wire445[(3'h5):(1'h1)])}));
            end
          reg456 <= $signed(((8'hab) ?
              (forvar448 <= $unsigned((8'hbb))) : $signed($signed(forvar452))));
          if ($signed((wire447[(3'h4):(2'h2)] << (wire446 ?
              wire445[(3'h5):(1'h0)] : $signed(((8'hb7) ? reg454 : wire445))))))
            begin
              reg457 = "taCWd4TEnh06R4o0k";
              reg458 <= wire444[(3'h7):(1'h0)];
            end
          else
            begin
              reg457 = $signed($signed($signed({$unsigned(wire446),
                  {forvar448}})));
              reg458 <= $signed((+(forvar448[(4'hd):(4'hd)] ?
                  wire446 : $signed(forvar452[(3'h4):(1'h0)]))));
              reg459 = "5MdKacuuBR";
              reg460 <= wire444;
              reg461 <= {$signed(reg458)};
            end
          reg462 <= ((forvar448 ?
                  $signed((|(7'h44))) : (((forvar452 - wire444) && (wire447 ?
                          reg460 : wire446)) ?
                      $unsigned({wire444}) : wire447[(3'h7):(3'h7)])) ?
              (~^reg450) : (^(wire444[(4'he):(3'h4)] | reg460)));
          reg463 <= (reg459[(3'h6):(2'h2)] ?
              $unsigned(({$signed(reg455)} ?
                  $unsigned((|forvar451)) : ((8'ha4) ?
                      $unsigned((8'hb1)) : (reg459 ?
                          wire443 : reg462)))) : reg458[(1'h1):(1'h0)]);
        end
      for (forvar464 = (1'h0); (forvar464 < (1'h0)); forvar464 = (forvar464 + (1'h1)))
        begin
          if (wire443[(3'h4):(2'h2)])
            begin
              reg465 <= $signed((((reg462[(3'h7):(3'h5)] ?
                  ((7'h42) + reg460) : reg462[(4'he):(4'hd)]) <= forvar449[(3'h4):(2'h3)]) < {$unsigned((wire443 ?
                      (8'hb0) : wire443)),
                  reg453}));
            end
          else
            begin
              reg465 = $signed($unsigned($unsigned($signed($signed(reg458)))));
            end
          for (forvar466 = (1'h0); (forvar466 < (2'h2)); forvar466 = (forvar466 + (1'h1)))
            begin
              reg467 <= ((7'h40) <<< ($unsigned($signed({(8'hab)})) ?
                  reg455 : $unsigned($signed(forvar452))));
            end
        end
      for (forvar468 = (1'h0); (forvar468 < (2'h2)); forvar468 = (forvar468 + (1'h1)))
        begin
          for (forvar469 = (1'h0); (forvar469 < (3'h4)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 = wire447;
              reg471 <= $unsigned(reg460[(2'h2):(1'h1)]);
              reg472 <= $unsigned(("VdRFZz4E" > {(((8'hb8) ?
                      reg460 : (7'h42)) <<< (wire443 ? reg461 : (8'ha3))),
                  wire447[(4'hd):(4'ha)]}));
              reg473 <= (reg458[(2'h2):(1'h0)] ?
                  $signed(reg470[(3'h5):(2'h2)]) : (^~reg462));
            end
          for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
            begin
              reg475 = "GDiY8uzz2sQu4T9WV";
              reg476 = reg450[(4'h9):(1'h1)];
              reg477 <= {(^reg465[(3'h4):(1'h0)])};
              reg478 = (&($unsigned("z") ? forvar452 : reg460));
            end
          for (forvar479 = (1'h0); (forvar479 < (1'h1)); forvar479 = (forvar479 + (1'h1)))
            begin
              reg480 <= {"btcQK1",
                  ($signed((&{reg460})) - $signed(reg472[(2'h2):(2'h2)]))};
            end
        end
      for (forvar481 = (1'h0); (forvar481 < (3'h4)); forvar481 = (forvar481 + (1'h1)))
        begin
          if ({$signed(((~^(&reg458)) >>> ((-reg477) ?
                  $unsigned(forvar466) : $unsigned((8'hb9)))))})
            begin
              reg482 = (reg463[(3'h4):(1'h0)] > (forvar474 - $unsigned(wire444)));
              reg483 = (8'hb8);
              reg484 = wire447;
            end
          else
            begin
              reg482 = $unsigned({(((wire446 ? reg472 : reg463) <<< (reg470 ?
                      (8'ha0) : wire444)) > {((8'hac) <<< reg484)}),
                  {$signed((wire443 < (8'hb0)))}});
              reg483 = $unsigned((^reg463[(3'h5):(1'h1)]));
            end
          if (reg472)
            begin
              reg485 = (^~(!$unsigned(((reg460 ^ reg457) <<< (reg478 <= reg463)))));
              reg486 <= (reg483 ?
                  ((|(|(reg458 ^ forvar448))) ?
                      forvar468[(3'h5):(2'h2)] : ($unsigned((reg457 ?
                          reg453 : (8'ha5))) ~^ reg467[(4'ha):(1'h1)])) : (((8'hb2) < reg461) ?
                      $unsigned(((wire445 ? (8'hb5) : reg457) ?
                          wire446[(3'h5):(1'h0)] : (&forvar479))) : reg472[(2'h2):(1'h0)]));
            end
          else
            begin
              reg485 = $unsigned(forvar481);
              reg486 <= reg482;
              reg487 <= "ZPPdTAv";
              reg488 <= $signed($signed((-($signed(reg470) ?
                  (-wire444) : (^forvar449)))));
              reg489 = reg475[(4'h8):(2'h3)];
            end
        end
    end
  assign wire490 = (wire443[(4'h9):(3'h6)] ?
                       $unsigned($signed(($signed(reg465) ?
                           {reg472} : (|(8'hb3))))) : ($unsigned(reg484[(4'h8):(1'h1)]) ?
                           $unsigned(forvar481) : {((|forvar449) == reg485),
                               $signed(reg454[(3'h4):(2'h3)])}));
  assign wire491 = ((reg489 ?
                           $unsigned(((forvar448 >>> (8'ha6)) ?
                               forvar481[(1'h1):(1'h0)] : reg467)) : ((+reg484[(2'h2):(1'h0)]) << forvar469)) ?
                       $signed(({{wire444},
                           $signed(reg462)} - $unsigned("6rqD"))) : "LHqxJcBsHzX");
  always
    @(posedge clk) begin
      for (forvar492 = (1'h0); (forvar492 < (2'h3)); forvar492 = (forvar492 + (1'h1)))
        begin
          for (forvar493 = (1'h0); (forvar493 < (1'h1)); forvar493 = (forvar493 + (1'h1)))
            begin
              reg494 <= $signed($unsigned(((wire444 != $signed(reg485)) ?
                  (8'hab) : forvar493[(2'h3):(1'h1)])));
            end
          reg495 <= $unsigned({(8'hab),
              $signed(((reg494 ? reg456 : wire490) ^ $unsigned(forvar452)))});
          for (forvar496 = (1'h0); (forvar496 < (3'h4)); forvar496 = (forvar496 + (1'h1)))
            begin
              reg497 = forvar448[(4'hb):(1'h0)];
              reg498 <= $signed(("f3dihrZf7TWlAP" >>> (($unsigned(reg459) ?
                      {reg457, (8'hb9)} : (wire446 > (8'hb2))) ?
                  reg461[(3'h5):(1'h1)] : {reg476})));
            end
          reg499 = wire491[(3'h6):(2'h2)];
          reg500 = (^$signed(forvar451[(1'h1):(1'h0)]));
        end
      reg501 = (reg472[(3'h4):(1'h1)] & forvar469[(4'ha):(3'h7)]);
      reg502 <= (((forvar468[(4'hd):(2'h3)] ?
          reg501 : $signed((forvar474 ? forvar493 : forvar492))) != (^((8'hb1) ?
          (|wire443) : {reg462,
              reg450}))) * $unsigned({($signed(reg486) + forvar492[(1'h1):(1'h1)]),
          (^~$unsigned(reg485))}));
    end
  assign wire503 = $signed((reg499 ^ $unsigned((+(-reg465)))));
  always
    @(posedge clk) begin
      reg504 <= (-($unsigned({(forvar464 ? reg470 : reg482),
          ((8'hb3) ? forvar452 : forvar452)}) - ({{reg457},
          wire443[(4'h8):(2'h2)]} != forvar479)));
      for (forvar505 = (1'h0); (forvar505 < (3'h4)); forvar505 = (forvar505 + (1'h1)))
        begin
          reg506 <= forvar452[(4'hd):(4'h9)];
          for (forvar507 = (1'h0); (forvar507 < (1'h1)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 = $signed((reg484 ?
                  {$unsigned(reg465)} : ($signed((-wire443)) <= (~$unsigned(forvar449)))));
              reg509 <= $unsigned($signed(reg461[(4'h8):(3'h4)]));
              reg510 = ((reg498[(2'h3):(1'h0)] || reg506[(3'h6):(2'h2)]) ?
                  (8'haf) : forvar481);
              reg511 <= (^~wire503);
            end
          reg512 <= wire490[(4'ha):(2'h3)];
        end
      reg513 <= reg450;
      for (forvar514 = (1'h0); (forvar514 < (1'h0)); forvar514 = (forvar514 + (1'h1)))
        begin
          if ($signed($signed(wire503)))
            begin
              reg515 <= forvar448;
            end
          else
            begin
              reg515 <= {((+forvar464[(3'h5):(2'h3)]) || $unsigned($unsigned((reg513 ?
                      forvar505 : reg455)))),
                  ($signed(reg453[(1'h0):(1'h0)]) ?
                      reg485[(1'h1):(1'h1)] : $signed((!$unsigned(reg463))))};
              reg516 <= ({$unsigned((~|(reg513 ?
                      forvar481 : reg465)))} >>> $unsigned(((~&reg500) && reg459)));
              reg517 = reg512[(4'hf):(4'hd)];
              reg518 = $signed(($unsigned($signed((reg494 ?
                      forvar493 : reg456))) ?
                  (8'hbb) : $signed((reg461 & reg500))));
            end
          for (forvar519 = (1'h0); (forvar519 < (3'h4)); forvar519 = (forvar519 + (1'h1)))
            begin
              reg520 = $signed({reg461[(2'h3):(1'h1)]});
              reg521 = (wire444 ?
                  reg467 : $signed($unsigned(({(8'ha9), reg456} - reg494))));
            end
          for (forvar522 = (1'h0); (forvar522 < (1'h0)); forvar522 = (forvar522 + (1'h1)))
            begin
              reg523 <= forvar469[(3'h5):(1'h1)];
              reg524 <= (-reg478);
            end
          if ((+$unsigned((($signed(reg523) ?
              $signed((8'ha7)) : reg520[(1'h0):(1'h0)]) ^~ (!"tA")))))
            begin
              reg525 <= $signed($signed(($unsigned((reg478 ?
                  reg473 : forvar464)) <<< (&(+wire447)))));
              reg526 <= reg498;
              reg527 <= $unsigned(reg520);
            end
          else
            begin
              reg525 <= ((~($unsigned(forvar481) - {$unsigned(reg506),
                  (reg495 == (8'h9f))})) >> reg483);
              reg526 <= ($unsigned(reg521[(3'h6):(1'h1)]) >> "0faTp");
              reg527 = ({reg484,
                  $unsigned($signed((reg504 & forvar492)))} && $signed($unsigned(reg477)));
            end
          for (forvar528 = (1'h0); (forvar528 < (1'h1)); forvar528 = (forvar528 + (1'h1)))
            begin
              reg529 <= (&$unsigned($unsigned(reg460)));
              reg530 = ((~&((|reg526) ?
                  {$unsigned(wire445),
                      $signed(reg500)} : reg518[(2'h2):(2'h2)])) << reg460);
              reg531 <= $signed($signed(((~&forvar505) != ($signed(reg504) ?
                  (forvar481 || reg498) : $unsigned(reg520)))));
            end
        end
      reg532 <= (~^(({{forvar468}} && reg465) << {($signed(reg531) ?
              $unsigned(reg471) : (reg459 < reg467))}));
    end
  always
    @(posedge clk) begin
      if ((({reg517[(2'h2):(2'h2)]} ?
              (((|reg501) >= (forvar505 ? (8'hab) : reg488)) ?
                  (8'ha3) : forvar514[(1'h1):(1'h1)]) : (($unsigned(reg512) ?
                      $signed(wire443) : $unsigned(reg532)) ?
                  reg516 : wire491[(1'h1):(1'h1)])) ?
          "f6k16xCZVYEg" : $signed((((forvar466 ? (7'h43) : reg480) ?
              (-reg524) : $signed((8'ha9))) ^ {{reg486}}))))
        begin
          for (forvar533 = (1'h0); (forvar533 < (2'h3)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 <= (^(reg521[(5'h11):(5'h11)] > ($unsigned($signed(reg489)) <<< $signed($unsigned((8'ha9))))));
              reg535 = $unsigned($signed((+wire503)));
            end
          if ((!forvar451[(2'h2):(1'h0)]))
            begin
              reg536 = reg488[(3'h7):(1'h0)];
              reg537 <= $signed(($signed((-$signed(forvar496))) <= forvar528));
              reg538 = $signed(wire445[(3'h5):(2'h3)]);
            end
          else
            begin
              reg536 <= {((reg453[(4'hd):(1'h1)] - (~&$signed(reg508))) ?
                      $unsigned(reg510) : reg523)};
              reg537 <= (reg450[(3'h7):(1'h1)] ?
                  $signed(forvar448) : (!$unsigned(reg537)));
              reg538 <= $unsigned($unsigned(forvar466[(2'h3):(1'h0)]));
              reg539 <= reg465;
            end
          for (forvar540 = (1'h0); (forvar540 < (1'h0)); forvar540 = (forvar540 + (1'h1)))
            begin
              reg541 <= reg518[(4'h8):(1'h1)];
              reg542 = (!(($signed(reg539) | {reg482[(1'h0):(1'h0)],
                  (&reg476)}) >>> reg461[(3'h4):(2'h3)]));
              reg543 = $signed(forvar449);
              reg544 <= "oI6aXFQ";
            end
          reg545 = reg456[(2'h2):(1'h1)];
          for (forvar546 = (1'h0); (forvar546 < (2'h3)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = ((^~(~|$unsigned({(8'h9e),
                  (8'hab)}))) << {((~^(forvar469 <<< reg531)) == (reg535 ?
                      (reg478 * (8'hb0)) : reg488[(1'h0):(1'h0)])),
                  (reg531 ?
                      (~$unsigned(reg472)) : $signed((wire446 ?
                          reg462 : (8'ha1))))});
            end
        end
      else
        begin
          for (forvar533 = (1'h0); (forvar533 < (2'h3)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 <= {reg485};
              reg535 <= (|(&(reg545[(4'hb):(4'h8)] ?
                  $unsigned((forvar469 ?
                      reg512 : wire490)) : (reg499 >>> "KusFB2m1rAy"))));
            end
          for (forvar536 = (1'h0); (forvar536 < (1'h1)); forvar536 = (forvar536 + (1'h1)))
            begin
              reg537 <= (-(reg454 ^~ {($signed((8'ha4)) ~^ (reg517 ~^ forvar496))}));
              reg538 <= $unsigned($signed($unsigned(reg516[(4'h8):(1'h1)])));
              reg539 = (reg484 != forvar474);
              reg540 <= reg459;
              reg541 = ((~|$unsigned((reg472 | $signed(reg454)))) ?
                  (reg540[(4'h8):(1'h1)] ?
                      $signed(reg470[(4'hd):(4'hc)]) : reg494[(2'h3):(2'h3)]) : $signed(reg494[(1'h0):(1'h0)]));
            end
          for (forvar542 = (1'h0); (forvar542 < (1'h0)); forvar542 = (forvar542 + (1'h1)))
            begin
              reg543 = ($unsigned($unsigned((!$unsigned(reg484)))) ?
                  (8'hb7) : ((reg467[(3'h6):(1'h0)] ?
                          (!reg508[(2'h2):(1'h1)]) : (reg508 ~^ $signed(reg525))) ?
                      (reg501[(2'h2):(1'h0)] ?
                          reg467[(1'h1):(1'h0)] : (^~"Bk")) : $unsigned({$unsigned(wire444),
                          (-forvar496)})));
            end
        end
    end
  assign wire548 = reg457[(4'h9):(3'h6)];
  always
    @(posedge clk) begin
      if ((forvar540 || $signed(reg453[(3'h6):(1'h1)])))
        begin
          for (forvar549 = (1'h0); (forvar549 < (2'h2)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= (reg461[(2'h3):(1'h0)] ?
                  $unsigned((!reg494)) : $signed((&$signed((reg484 || reg516)))));
              reg551 = (reg459 ?
                  (forvar452 ?
                      $signed(forvar546[(1'h1):(1'h1)]) : {reg455}) : $signed($signed($signed(forvar479))));
            end
          for (forvar552 = (1'h0); (forvar552 < (1'h1)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 <= ($unsigned($unsigned($signed((forvar536 ^ reg488)))) ?
                  (reg499 ?
                      (|reg550) : (forvar507 ~^ reg489[(2'h2):(1'h1)])) : reg544);
              reg554 <= reg536[(3'h4):(2'h3)];
              reg555 <= (reg551 - $signed({$signed(wire447)}));
            end
        end
      else
        begin
          for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 = $signed($signed($signed(($unsigned(reg535) ^~ forvar449[(2'h3):(2'h2)]))));
            end
          for (forvar551 = (1'h0); (forvar551 < (3'h4)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 <= ($signed(reg450[(2'h2):(1'h1)]) >= forvar451);
              reg553 = ($signed(wire447) >> forvar449);
            end
          for (forvar554 = (1'h0); (forvar554 < (1'h1)); forvar554 = (forvar554 + (1'h1)))
            begin
              reg555 <= $unsigned($unsigned(reg544[(1'h1):(1'h0)]));
            end
        end
      for (forvar556 = (1'h0); (forvar556 < (1'h0)); forvar556 = (forvar556 + (1'h1)))
        begin
          for (forvar557 = (1'h0); (forvar557 < (1'h1)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 <= forvar552;
            end
          reg559 = reg504[(3'h4):(2'h3)];
          for (forvar560 = (1'h0); (forvar560 < (3'h4)); forvar560 = (forvar560 + (1'h1)))
            begin
              reg561 <= ($signed((~^$signed((|reg559)))) <<< $unsigned((((^reg516) ?
                      forvar551 : {wire445}) ?
                  $signed($unsigned(forvar496)) : reg455[(1'h1):(1'h0)])));
            end
          reg562 = $signed((({$signed((8'hbb)),
              reg553} ^~ forvar554) < (^~forvar533[(3'h5):(2'h3)])));
          reg563 = forvar552;
        end
      reg564 <= (reg540 || reg475);
    end
  assign wire565 = (reg462[(3'h5):(3'h5)] <<< forvar551[(4'h8):(4'h8)]);
  always
    @(posedge clk) begin
      reg566 = $unsigned((reg512[(1'h0):(1'h0)] ?
          "FF8DXI0" : ((reg547[(1'h0):(1'h0)] ?
              (reg535 ?
                  reg459 : reg460) : $unsigned(reg488)) ^ $signed(reg454))));
      reg567 <= ((~&$signed({(forvar505 ^~ reg483)})) ~^ reg525[(2'h3):(1'h1)]);
      for (forvar568 = (1'h0); (forvar568 < (2'h3)); forvar568 = (forvar568 + (1'h1)))
        begin
          reg569 = reg470[(1'h1):(1'h1)];
          reg570 = reg498[(2'h2):(2'h2)];
          for (forvar571 = (1'h0); (forvar571 < (3'h4)); forvar571 = (forvar571 + (1'h1)))
            begin
              reg572 = (^~$unsigned($signed((&(~&forvar549)))));
              reg573 <= reg530;
              reg574 <= $signed($unsigned($unsigned(reg494[(1'h1):(1'h0)])));
            end
          for (forvar575 = (1'h0); (forvar575 < (3'h4)); forvar575 = (forvar575 + (1'h1)))
            begin
              reg576 <= $unsigned(($signed($signed("")) * reg489[(2'h2):(2'h2)]));
              reg577 <= "KVZn2O11is2aPzVmzn";
              reg578 <= {wire443[(4'h9):(4'h8)],
                  {$unsigned((-((8'hac) ? reg473 : forvar505))),
                      $unsigned(forvar542[(2'h2):(2'h2)])}};
            end
          for (forvar579 = (1'h0); (forvar579 < (2'h3)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 = $signed($signed(forvar514[(5'h11):(3'h7)]));
            end
        end
      reg581 <= reg580[(3'h7):(1'h1)];
      for (forvar582 = (1'h0); (forvar582 < (2'h2)); forvar582 = (forvar582 + (1'h1)))
        begin
          reg583 <= $signed(((|(~&(reg526 ?
              reg526 : wire444))) && {$signed((|forvar493)),
              "VHXscqm5uhNQqH1"}));
          reg584 <= reg539[(2'h3):(2'h3)];
          reg585 = (~&$signed(reg558[(4'h9):(3'h7)]));
          reg586 <= $unsigned((|$signed($unsigned(reg470))));
        end
    end
  always
    @(posedge clk) begin
      reg587 = forvar481;
      if (reg515[(4'h8):(3'h5)])
        begin
          for (forvar588 = (1'h0); (forvar588 < (1'h0)); forvar588 = (forvar588 + (1'h1)))
            begin
              reg589 = forvar560;
              reg590 = reg450[(1'h1):(1'h0)];
              reg591 <= "pHQCMbfcEVGgvo";
              reg592 <= (&reg450[(4'h9):(3'h4)]);
            end
          for (forvar593 = (1'h0); (forvar593 < (2'h3)); forvar593 = (forvar593 + (1'h1)))
            begin
              reg594 <= (((&reg501[(3'h4):(3'h4)]) & {(~&(forvar479 | reg473))}) && (&$unsigned(((reg461 - reg517) < reg535))));
            end
        end
      else
        begin
          reg588 = (&(reg482 ? reg572[(3'h4):(3'h4)] : reg532));
          for (forvar589 = (1'h0); (forvar589 < (2'h3)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 <= (reg572 & (({(!(8'hbd)), {(8'ha8), (8'hbc)}} ?
                  $unsigned(reg525) : reg499) | reg460));
              reg591 <= {$signed({($signed(reg566) < $signed(reg472))}),
                  (reg534[(4'he):(4'hc)] ?
                      $unsigned((+(^~reg542))) : (reg453 ~^ (8'hb4)))};
              reg592 <= {reg537};
            end
        end
    end
  assign wire595 = (reg550[(4'h8):(4'h8)] && $unsigned($signed((^~{reg544}))));
  always
    @(posedge clk) begin
      if (reg559)
        begin
          for (forvar596 = (1'h0); (forvar596 < (1'h0)); forvar596 = (forvar596 + (1'h1)))
            begin
              reg597 <= wire565[(2'h2):(1'h0)];
            end
          for (forvar598 = (1'h0); (forvar598 < (2'h3)); forvar598 = (forvar598 + (1'h1)))
            begin
              reg599 <= $signed((+(reg587 ?
                  $signed($signed(reg454)) : (reg580 ?
                      (forvar596 ? reg450 : (8'ha5)) : {(8'hb5)}))));
              reg600 <= ($signed(reg518[(1'h0):(1'h0)]) | $unsigned(forvar519[(4'hd):(3'h5)]));
              reg601 <= reg457[(2'h3):(1'h1)];
              reg602 = {(~($signed($signed(forvar452)) ?
                      $unsigned(reg497[(2'h2):(1'h0)]) : ((reg495 || (7'h41)) ?
                          {reg471} : $signed(forvar528)))),
                  reg498};
            end
        end
      else
        begin
          reg596 = $signed({reg494[(1'h1):(1'h0)]});
          reg597 <= (reg502[(4'hb):(4'ha)] ^ reg450);
          reg598 <= (wire491 >>> $signed($unsigned(forvar593)));
          if ((^~$unsigned($unsigned(reg554))))
            begin
              reg599 = ((8'hae) ?
                  {($unsigned($unsigned(forvar579)) ?
                          $unsigned(forvar474) : ((reg551 ? reg600 : (8'hb0)) ?
                              {reg591} : forvar542)),
                      $signed($signed(forvar552))} : (reg485[(3'h5):(1'h0)] >>> ($unsigned((forvar493 - reg520)) ?
                      reg563[(4'hb):(4'h9)] : $unsigned((reg453 ?
                          (8'hbe) : forvar557)))));
              reg600 = {reg488[(4'h8):(3'h4)],
                  $signed((~^$signed((&forvar493))))};
              reg601 = {(~(^~((wire490 ? forvar582 : reg592) ?
                      (wire444 != (8'hb0)) : (|reg598)))),
                  reg564};
              reg602 = (~|$unsigned("Froz5DKI"));
              reg603 = {({$signed((~(7'h44)))} <<< $signed($unsigned($signed(forvar596))))};
            end
          else
            begin
              reg599 = forvar507;
              reg600 = forvar579;
              reg601 = $signed(forvar579[(1'h1):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar604 = (1'h0); (forvar604 < (3'h4)); forvar604 = (forvar604 + (1'h1)))
        begin
          reg605 = (!(reg594[(4'h9):(1'h0)] ?
              {$unsigned($unsigned(reg577)),
                  ($signed(reg498) ?
                      (forvar474 ~^ reg599) : forvar604)} : $unsigned($unsigned(forvar554))));
          reg606 <= wire565[(2'h2):(1'h0)];
          if ($unsigned((8'hba)))
            begin
              reg607 <= (reg502[(3'h5):(1'h0)] * forvar474);
              reg608 <= forvar493;
            end
          else
            begin
              reg607 = ($signed(reg550) ?
                  $unsigned((~&reg470)) : $unsigned(($signed(reg510[(1'h1):(1'h0)]) ?
                      "5NMpdSdPCrAKIm3MY9Ls" : $unsigned($unsigned(reg596)))));
              reg608 <= $unsigned({$unsigned((~$signed(forvar589))),
                  ($signed((^(7'h42))) ?
                      wire443[(1'h0):(1'h0)] : $unsigned($unsigned(forvar589)))});
              reg609 = (^(|($unsigned($signed(reg541)) >= ($signed(wire503) ?
                  reg463 : $signed(reg555)))));
              reg610 <= (("o" ?
                  (8'h9c) : (^($signed(reg526) * reg597[(2'h2):(2'h2)]))) << (7'h42));
              reg611 <= $unsigned((^$signed($signed({(8'h9e), (8'haa)}))));
            end
          for (forvar612 = (1'h0); (forvar612 < (1'h0)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 <= "byr";
              reg614 <= forvar557[(3'h5):(3'h5)];
              reg615 <= ($unsigned(reg508) ?
                  ($signed(reg605) ?
                      ($signed(((8'ha6) ? forvar528 : forvar568)) ?
                          $signed($unsigned(reg462)) : ($unsigned((8'hbf)) ?
                              (~|forvar546) : $signed(reg450))) : (reg538 ^ (7'h41))) : $signed(reg486));
              reg616 <= (reg482[(4'ha):(3'h4)] * $signed(($unsigned((reg506 > reg607)) ?
                  ({forvar449} ^~ forvar449[(2'h3):(1'h0)]) : reg455)));
              reg617 = reg537;
            end
        end
      for (forvar618 = (1'h0); (forvar618 < (3'h4)); forvar618 = (forvar618 + (1'h1)))
        begin
          reg619 <= reg545[(2'h2):(1'h1)];
          reg620 = forvar536;
          for (forvar621 = (1'h0); (forvar621 < (2'h3)); forvar621 = (forvar621 + (1'h1)))
            begin
              reg622 <= reg524[(3'h5):(1'h1)];
            end
          reg623 <= $unsigned(($signed($signed($unsigned((8'h9f)))) >>> forvar507[(4'hf):(4'h8)]));
          reg624 = $unsigned(reg524[(2'h2):(1'h1)]);
        end
      reg625 <= reg601[(3'h4):(1'h0)];
      reg626 = {$unsigned("TRPA4eHaWHVIFGcGx7"),
          ({(~^(~forvar449)), $signed(forvar618)} ?
              (reg489[(2'h2):(1'h1)] ?
                  "hkd" : ((!(8'ha9)) ?
                      (reg570 >>> forvar519) : (reg520 ?
                          forvar468 : reg534))) : reg623[(4'ha):(1'h1)])};
      for (forvar627 = (1'h0); (forvar627 < (1'h0)); forvar627 = (forvar627 + (1'h1)))
        begin
          if ((reg544 - $signed($unsigned($signed((reg538 ?
              reg457 : reg512))))))
            begin
              reg628 <= ((^$unsigned($signed(((8'hae) ? reg495 : forvar621)))) ?
                  $signed(($signed($signed((8'ha7))) ?
                      ((reg554 ?
                          reg460 : reg525) || $signed(reg609)) : reg603[(1'h1):(1'h1)])) : $signed(($signed((reg477 ?
                      (8'ha8) : reg543)) >> {(reg504 != forvar451),
                      forvar528[(1'h0):(1'h0)]})));
              reg629 <= $signed($unsigned(reg459));
              reg630 = (((forvar598[(4'hb):(4'hb)] ?
                      reg624 : (forvar575 ?
                          $unsigned(forvar588) : (&forvar505))) > ((+$unsigned((8'hb3))) ?
                      (~^$unsigned(reg456)) : $unsigned(wire443))) ?
                  reg622 : $signed($signed($signed((^reg545)))));
            end
          else
            begin
              reg628 = ($unsigned($signed(({reg477, reg613} ?
                  (reg527 >= reg569) : (forvar481 ?
                      reg551 : reg553)))) != (reg536[(5'h14):(4'hc)] ?
                  $unsigned(((~reg562) << {reg543})) : {((reg535 != forvar533) || reg525),
                      {((8'hac) ? forvar519 : reg482),
                          (reg480 ? forvar448 : reg570)}}));
              reg629 = $signed({(|($unsigned(reg517) ?
                      (reg563 ? reg581 : reg551) : (8'h9f))),
                  (reg559[(2'h2):(2'h2)] ? $unsigned(reg613) : forvar604)});
              reg630 <= $signed(forvar549[(4'hf):(4'hb)]);
            end
          for (forvar631 = (1'h0); (forvar631 < (1'h1)); forvar631 = (forvar631 + (1'h1)))
            begin
              reg632 <= reg542;
              reg633 = (~&reg524);
              reg634 = reg547;
              reg635 <= (reg620 < {(~&reg534[(3'h6):(3'h4)])});
            end
          for (forvar636 = (1'h0); (forvar636 < (2'h3)); forvar636 = (forvar636 + (1'h1)))
            begin
              reg637 <= $unsigned((+$signed($signed((reg578 ?
                  reg457 : forvar546)))));
              reg638 <= (^{$unsigned("p6hueFWk9hTNz1SZZaq"), $signed(reg537)});
              reg639 <= (8'ha1);
              reg640 <= ({(~&{$unsigned(forvar514), $unsigned(reg504)}),
                  reg606[(1'h0):(1'h0)]} << $signed(({reg523[(3'h7):(2'h2)],
                      (8'ha4)} ?
                  (-reg639[(2'h3):(2'h3)]) : "QL4GhXG")));
            end
        end
    end
  assign wire641 = forvar546[(1'h1):(1'h0)];
endmodule
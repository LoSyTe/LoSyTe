(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param679 = ({(~(~|(~^(8'hb0)))), (((|(8'had)) + ((8'hb0) && (8'hb7))) >= (~^((8'ha4) ? (8'haf) : (8'h9f))))} - ({({(7'h40), (8'hb9)} ? ((8'hb6) ? (8'h9e) : (8'h9e)) : ((8'hb9) || (8'hab))), ({(8'ha8)} ? ((8'hb8) ? (8'hb2) : (8'h9c)) : {(7'h44), (8'hb3)})} ? ((+((8'ha7) ? (8'hb3) : (8'h9e))) ? {((8'hb7) ^~ (8'hb9)), ((7'h41) ? (8'ha6) : (8'hbb))} : {((7'h42) < (8'ha1)), {(7'h41)}}) : (|(~&((8'ha2) ? (8'hbe) : (8'h9c))))))
, parameter param680 = ({(((param679 ? (8'h9f) : param679) ^ {param679, (8'ha5)}) ? (~^{param679, (8'hab)}) : ((param679 >= param679) ? (param679 ? param679 : param679) : (param679 ? param679 : param679)))} || ((param679 <= (param679 == (param679 ? param679 : param679))) ? {param679, param679} : (!param679))) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h9d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire4;
  input wire signed [(3'h4):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire2;
  input wire [(4'he):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire0;
  wire [(4'hb):(1'h0)] wire677;
  wire signed [(5'h13):(1'h0)] wire676;
  reg signed [(5'h15):(1'h0)] reg675 = (1'h0);
  reg [(5'h15):(1'h0)] forvar674 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire605;
  reg signed [(4'hc):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg603 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire602;
  reg signed [(2'h3):(1'h0)] reg601 = (1'h0);
  reg signed [(4'he):(1'h0)] reg600 = (1'h0);
  reg [(3'h5):(1'h0)] reg599 = (1'h0);
  reg [(3'h4):(1'h0)] forvar598 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar597 = (1'h0);
  reg [(4'hb):(1'h0)] reg596 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar595 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg594 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg593 = (1'h0);
  reg [(5'h12):(1'h0)] reg592 = (1'h0);
  reg [(4'hf):(1'h0)] forvar591 = (1'h0);
  reg [(5'h15):(1'h0)] reg590 = (1'h0);
  reg [(5'h12):(1'h0)] reg589 = (1'h0);
  reg [(4'hb):(1'h0)] reg588 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg587 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg585 = (1'h0);
  reg [(4'hf):(1'h0)] forvar584 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar583 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg581 = (1'h0);
  reg [(4'hc):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar579 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg578 = (1'h0);
  reg [(4'hf):(1'h0)] reg577 = (1'h0);
  reg [(3'h7):(1'h0)] reg576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg575 = (1'h0);
  reg [(5'h12):(1'h0)] reg574 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar573 = (1'h0);
  reg [(5'h13):(1'h0)] reg572 = (1'h0);
  reg [(4'he):(1'h0)] forvar571 = (1'h0);
  reg [(3'h4):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg561 = (1'h0);
  reg [(4'hb):(1'h0)] reg557 = (1'h0);
  reg [(5'h11):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar553 = (1'h0);
  reg [(3'h6):(1'h0)] reg569 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg568 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg566 = (1'h0);
  reg [(2'h2):(1'h0)] reg565 = (1'h0);
  reg [(3'h7):(1'h0)] forvar564 = (1'h0);
  reg [(4'hb):(1'h0)] reg563 = (1'h0);
  reg [(5'h15):(1'h0)] reg562 = (1'h0);
  reg [(5'h15):(1'h0)] forvar561 = (1'h0);
  reg [(5'h13):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg559 = (1'h0);
  reg [(2'h2):(1'h0)] reg558 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar557 = (1'h0);
  reg [(5'h11):(1'h0)] reg556 = (1'h0);
  reg signed [(4'he):(1'h0)] reg555 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar554 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg553 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire552;
  wire [(3'h4):(1'h0)] wire551;
  reg signed [(4'he):(1'h0)] reg550 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg549 = (1'h0);
  reg [(4'he):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg547 = (1'h0);
  reg [(5'h15):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg545 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg544 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg543 = (1'h0);
  reg [(2'h3):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar541 = (1'h0);
  reg [(5'h11):(1'h0)] reg540 = (1'h0);
  reg [(5'h15):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar538 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg537 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar536 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg535 = (1'h0);
  reg [(5'h10):(1'h0)] reg534 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg533 = (1'h0);
  reg [(5'h10):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar531 = (1'h0);
  reg [(4'hf):(1'h0)] reg530 = (1'h0);
  reg [(4'hf):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg528 = (1'h0);
  reg [(4'hc):(1'h0)] reg527 = (1'h0);
  reg [(4'h8):(1'h0)] reg526 = (1'h0);
  reg [(3'h4):(1'h0)] reg525 = (1'h0);
  reg [(4'h8):(1'h0)] reg524 = (1'h0);
  reg [(5'h15):(1'h0)] forvar523 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg522 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg521 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg520 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg519 = (1'h0);
  reg [(3'h5):(1'h0)] reg518 = (1'h0);
  reg [(4'ha):(1'h0)] forvar517 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar516 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg515 = (1'h0);
  reg [(4'h8):(1'h0)] forvar514 = (1'h0);
  reg [(4'h9):(1'h0)] reg513 = (1'h0);
  reg [(5'h14):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg511 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg510 = (1'h0);
  reg [(2'h2):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg508 = (1'h0);
  reg [(3'h5):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar506 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg505 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg504 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg503 = (1'h0);
  reg [(2'h3):(1'h0)] forvar502 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg501 = (1'h0);
  reg [(5'h14):(1'h0)] forvar500 = (1'h0);
  reg [(5'h11):(1'h0)] reg499 = (1'h0);
  reg [(2'h3):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg497 = (1'h0);
  reg [(4'he):(1'h0)] reg496 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg495 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg494 = (1'h0);
  reg [(3'h5):(1'h0)] reg493 = (1'h0);
  reg [(5'h14):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar491 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar490 = (1'h0);
  reg [(3'h4):(1'h0)] reg489 = (1'h0);
  wire [(2'h2):(1'h0)] wire60;
  reg signed [(5'h13):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg12 = (1'h0);
  reg [(5'h14):(1'h0)] reg11 = (1'h0);
  reg [(3'h6):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg9 = (1'h0);
  reg [(3'h6):(1'h0)] reg8 = (1'h0);
  reg [(4'hd):(1'h0)] reg7 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire487;
  reg signed [(5'h10):(1'h0)] reg607 = (1'h0);
  reg [(4'hc):(1'h0)] forvar608 = (1'h0);
  reg [(4'hd):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar610 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar611 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg613 = (1'h0);
  reg [(4'hd):(1'h0)] forvar614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg615 = (1'h0);
  reg [(5'h15):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar618 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg619 = (1'h0);
  reg [(3'h7):(1'h0)] reg620 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg622 = (1'h0);
  reg [(3'h4):(1'h0)] forvar623 = (1'h0);
  reg [(3'h7):(1'h0)] reg624 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg627 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar629 = (1'h0);
  reg [(5'h12):(1'h0)] reg630 = (1'h0);
  reg [(4'he):(1'h0)] reg631 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire632;
  reg signed [(5'h14):(1'h0)] forvar633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg634 = (1'h0);
  reg [(5'h15):(1'h0)] reg635 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar637 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg638 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg639 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg641 = (1'h0);
  reg [(2'h3):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg643 = (1'h0);
  reg [(5'h14):(1'h0)] reg644 = (1'h0);
  reg [(4'hb):(1'h0)] reg645 = (1'h0);
  reg [(3'h7):(1'h0)] forvar646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg647 = (1'h0);
  reg [(4'he):(1'h0)] reg648 = (1'h0);
  reg [(5'h10):(1'h0)] reg649 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg633 = (1'h0);
  reg signed [(4'he):(1'h0)] reg651 = (1'h0);
  reg [(5'h11):(1'h0)] forvar652 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar653 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg654 = (1'h0);
  reg [(5'h12):(1'h0)] reg655 = (1'h0);
  reg [(2'h3):(1'h0)] reg656 = (1'h0);
  reg [(5'h14):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg658 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar659 = (1'h0);
  reg [(4'hb):(1'h0)] reg660 = (1'h0);
  reg [(4'hf):(1'h0)] reg661 = (1'h0);
  reg [(5'h13):(1'h0)] forvar662 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg664 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg665 = (1'h0);
  reg [(5'h12):(1'h0)] reg666 = (1'h0);
  reg [(5'h12):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar669 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg670 = (1'h0);
  reg [(4'h9):(1'h0)] reg662 = (1'h0);
  reg [(3'h6):(1'h0)] forvar663 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar665 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire671;
  wire [(5'h11):(1'h0)] wire672;
  assign y = {wire677,
                 wire676,
                 reg675,
                 forvar674,
                 wire605,
                 reg604,
                 reg603,
                 wire602,
                 reg601,
                 reg600,
                 reg599,
                 forvar598,
                 forvar597,
                 reg596,
                 forvar595,
                 reg594,
                 reg593,
                 reg592,
                 forvar591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 forvar584,
                 forvar583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 reg572,
                 forvar571,
                 reg570,
                 reg561,
                 reg557,
                 reg554,
                 forvar553,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 forvar564,
                 reg563,
                 reg562,
                 forvar561,
                 reg560,
                 reg559,
                 reg558,
                 forvar557,
                 reg556,
                 reg555,
                 forvar554,
                 reg553,
                 wire552,
                 wire551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 forvar541,
                 reg540,
                 reg539,
                 forvar538,
                 reg537,
                 forvar536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 forvar523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 forvar517,
                 forvar516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 forvar506,
                 reg505,
                 reg504,
                 reg503,
                 forvar502,
                 reg501,
                 forvar500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 forvar491,
                 forvar490,
                 reg489,
                 wire60,
                 reg6,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 forvar6,
                 reg5,
                 wire487,
                 reg607,
                 forvar608,
                 reg609,
                 forvar610,
                 forvar611,
                 reg612,
                 reg613,
                 forvar614,
                 reg615,
                 reg616,
                 reg617,
                 forvar618,
                 reg619,
                 reg620,
                 reg621,
                 reg622,
                 forvar623,
                 reg624,
                 reg625,
                 reg626,
                 reg627,
                 reg628,
                 forvar629,
                 reg630,
                 reg631,
                 wire632,
                 forvar633,
                 reg634,
                 reg635,
                 reg636,
                 forvar637,
                 reg638,
                 reg639,
                 forvar640,
                 reg641,
                 reg642,
                 reg643,
                 reg644,
                 reg645,
                 forvar646,
                 reg647,
                 reg648,
                 reg649,
                 reg650,
                 reg633,
                 reg651,
                 forvar652,
                 forvar653,
                 reg654,
                 reg655,
                 reg656,
                 reg657,
                 reg658,
                 forvar659,
                 reg660,
                 reg661,
                 forvar662,
                 reg663,
                 reg664,
                 reg665,
                 reg666,
                 reg667,
                 reg668,
                 forvar669,
                 reg670,
                 reg662,
                 forvar663,
                 forvar665,
                 wire671,
                 wire672,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire2[(1'h0):(1'h0)])
        begin
          reg5 <= (7'h42);
          for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 <= (7'h42);
              reg8 <= ((~|$signed($signed(wire3[(2'h3):(1'h1)]))) != $signed(reg7[(2'h2):(1'h1)]));
              reg9 <= wire4[(2'h3):(1'h1)];
              reg10 <= ({(8'h9d),
                  (^forvar6[(3'h4):(2'h3)])} >> (wire1[(3'h6):(3'h4)] ?
                  $unsigned(((wire1 || (8'hb7)) ^ wire3[(1'h0):(1'h0)])) : wire2[(2'h3):(2'h2)]));
              reg11 = $unsigned((&(&$unsigned({reg10}))));
            end
          reg12 <= ((forvar6[(4'hb):(1'h1)] && (&wire2[(3'h7):(3'h5)])) >>> ($unsigned(($unsigned(wire0) && $signed(reg8))) ?
              (wire1[(3'h6):(3'h4)] < wire1) : $signed($unsigned((reg10 >> reg5)))));
          reg13 <= $signed($unsigned((!$signed(((8'ha2) > wire3)))));
          reg14 <= {$signed((((reg12 ? reg8 : (8'ha4)) ?
                      forvar6[(4'hd):(3'h7)] : forvar6) ?
                  forvar6[(2'h2):(2'h2)] : $unsigned($unsigned(reg8)))),
              (!(~|$signed((7'h43))))};
        end
      else
        begin
          reg5 = {wire3[(1'h0):(1'h0)]};
          reg6 <= $unsigned((forvar6 ?
              ("KCPiaEMxJ" ?
                  wire0 : ((reg11 ?
                      wire2 : wire4) ~^ $unsigned(wire4))) : (~&(~&((8'h9f) ?
                  reg5 : wire4)))));
        end
    end
  module15 modinst61 (wire60, clk, wire2, reg9, reg14, reg12, reg5);
  module62 modinst488 (wire487, clk, wire2, reg7, wire1, wire0, forvar6);
  always
    @(posedge clk) begin
      reg489 <= $unsigned(($signed((-wire4)) >>> (8'hb9)));
      for (forvar490 = (1'h0); (forvar490 < (1'h0)); forvar490 = (forvar490 + (1'h1)))
        begin
          for (forvar491 = (1'h0); (forvar491 < (2'h3)); forvar491 = (forvar491 + (1'h1)))
            begin
              reg492 = $signed(reg6[(4'he):(4'h9)]);
              reg493 <= $unsigned($signed({(reg8 ?
                      $signed((8'h9c)) : {(8'ha7), reg14}),
                  $unsigned($signed(forvar491))}));
              reg494 = (!(~^$unsigned(($signed(reg13) ?
                  (~&(8'hbc)) : (reg13 ? reg10 : wire4)))));
              reg495 <= $signed(reg11[(1'h0):(1'h0)]);
              reg496 <= (8'hbb);
            end
          reg497 <= (((((^reg495) ? (-reg8) : (forvar6 ^ reg13)) ?
              {{reg14}, (reg6 >> reg11)} : $unsigned((reg13 ?
                  reg9 : (8'h9e)))) >> reg495) ^~ wire60[(2'h2):(1'h1)]);
        end
      reg498 <= ((({(wire0 || reg7)} ^ $signed(reg493[(2'h3):(2'h3)])) ?
          (wire0 ?
              (~wire1[(4'h8):(4'h8)]) : reg11) : (8'h9f)) >= ($signed(((reg492 ?
              reg5 : reg6) ?
          forvar490[(1'h1):(1'h1)] : (~|wire3))) == ({((8'ha8) | reg494),
              (reg13 ? wire2 : reg5)} ?
          wire2[(3'h6):(1'h0)] : ((&(8'hbd)) ~^ wire60))));
      reg499 <= $signed(("3pBlJ98Iaug" ^ wire3[(1'h0):(1'h0)]));
      for (forvar500 = (1'h0); (forvar500 < (2'h3)); forvar500 = (forvar500 + (1'h1)))
        begin
          reg501 = (((reg11 & $unsigned((reg6 ? reg499 : forvar6))) && reg10) ?
              $unsigned($signed((8'h9c))) : $signed(reg11));
          for (forvar502 = (1'h0); (forvar502 < (3'h4)); forvar502 = (forvar502 + (1'h1)))
            begin
              reg503 <= (&(8'ha7));
              reg504 = reg9;
              reg505 <= {$signed((~|$signed((+reg497))))};
            end
          for (forvar506 = (1'h0); (forvar506 < (2'h2)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 <= (8'ha3);
              reg508 = $unsigned((-(|{(reg503 - (8'hb8)), {wire2, reg7}})));
              reg509 = $unsigned((!$unsigned(((forvar502 ?
                  (7'h42) : wire60) ^~ reg499[(4'hc):(3'h7)]))));
              reg510 = (^(forvar502 ?
                  $signed(wire60) : ($unsigned({reg503}) ?
                      ((reg504 && wire1) | wire487) : reg503)));
              reg511 = (((reg7[(4'hb):(1'h0)] ?
                      reg13 : reg501[(4'hd):(4'ha)]) >> ((wire3[(2'h2):(1'h1)] <= ((8'hb8) >> reg505)) ?
                      reg8 : $unsigned((~&reg9)))) ?
                  $signed((reg12[(4'ha):(4'h8)] ?
                      reg504 : (~|((7'h40) & forvar500)))) : (~^(8'ha6)));
            end
          reg512 = ($unsigned(({$unsigned(forvar506)} ?
              reg499[(2'h3):(2'h2)] : reg498)) ^~ (~$unsigned($signed((^~reg510)))));
          reg513 <= ((&(~$unsigned((forvar6 ? (8'hb6) : forvar502)))) ?
              reg5 : reg499);
        end
    end
  always
    @(posedge clk) begin
      for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
        begin
          reg515 <= reg14;
        end
      for (forvar516 = (1'h0); (forvar516 < (3'h4)); forvar516 = (forvar516 + (1'h1)))
        begin
          for (forvar517 = (1'h0); (forvar517 < (1'h0)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 = (8'ha5);
              reg519 = $unsigned($signed("8MpC083g8lZa"));
              reg520 <= {reg14[(3'h4):(1'h0)]};
              reg521 = reg493;
            end
          reg522 <= reg495[(1'h0):(1'h0)];
          for (forvar523 = (1'h0); (forvar523 < (3'h4)); forvar523 = (forvar523 + (1'h1)))
            begin
              reg524 <= reg520;
              reg525 <= (reg505 ?
                  {(~^(reg503[(2'h2):(1'h0)] << $signed(reg507)))} : ($unsigned(reg497[(4'he):(3'h7)]) ?
                      $signed((~|(forvar502 + reg493))) : reg511));
              reg526 = (~^(($signed(wire2[(4'hb):(4'hb)]) != (reg525[(1'h0):(1'h0)] ?
                  (reg497 & wire487) : $signed(reg6))) == (("ZrfLtow5LzSpAeReRXZu" > $signed(reg520)) ?
                  {(wire0 ? (8'hae) : (8'hb2)), {reg519, reg505}} : (~|(reg8 ?
                      wire4 : reg493)))));
              reg527 = reg497;
              reg528 = forvar502[(2'h2):(1'h1)];
            end
          if (({$unsigned($unsigned({reg494}))} > $signed((wire0 ?
              $unsigned(reg521) : $unsigned((^~wire2))))))
            begin
              reg529 = "bGHtQY";
              reg530 <= (~&((~|reg497[(4'he):(3'h6)]) ?
                  ((~|reg509[(2'h2):(2'h2)]) ?
                      $unsigned((reg504 ?
                          reg528 : reg529)) : reg511) : (&(!reg526))));
            end
          else
            begin
              reg529 = (&reg518);
              reg530 = {"N6RRYgRGflcaS7El", reg513[(1'h0):(1'h0)]};
            end
          for (forvar531 = (1'h0); (forvar531 < (2'h2)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 = (^~forvar523[(5'h11):(2'h3)]);
              reg533 = $signed({$unsigned(((~|reg497) ?
                      $unsigned(reg530) : $unsigned(wire1))),
                  (|reg494[(2'h3):(2'h2)])});
              reg534 = reg505;
              reg535 <= (~|$signed(reg520));
            end
        end
      for (forvar536 = (1'h0); (forvar536 < (2'h3)); forvar536 = (forvar536 + (1'h1)))
        begin
          reg537 = (wire487[(3'h5):(1'h0)] ?
              $signed((-reg492[(2'h2):(2'h2)])) : (7'h41));
        end
      for (forvar538 = (1'h0); (forvar538 < (2'h2)); forvar538 = (forvar538 + (1'h1)))
        begin
          reg539 = $signed((forvar531 > (((reg495 || (7'h42)) ?
              (reg494 - (8'hb5)) : (8'hb2)) & ({reg527, reg496} ?
              $signed(forvar506) : {wire0, (8'hab)}))));
          reg540 = {forvar6[(3'h5):(1'h0)]};
          for (forvar541 = (1'h0); (forvar541 < (1'h0)); forvar541 = (forvar541 + (1'h1)))
            begin
              reg542 = (reg7 ~^ (^~(^forvar536)));
              reg543 <= "2nG";
              reg544 = $signed(reg505[(2'h3):(2'h2)]);
              reg545 <= reg522[(3'h6):(3'h4)];
            end
          if (reg543[(3'h4):(1'h0)])
            begin
              reg546 = (forvar500[(5'h12):(5'h12)] ^~ reg527[(2'h3):(1'h0)]);
              reg547 = wire1[(3'h5):(1'h0)];
              reg548 <= {"wLSy", $unsigned(reg505[(3'h6):(2'h3)])};
              reg549 = $unsigned((($signed({reg498, reg11}) ?
                      ($signed(reg503) > reg526) : reg526[(2'h2):(1'h1)]) ?
                  "RF9F63ba" : $unsigned(forvar516)));
              reg550 = wire4[(1'h0):(1'h0)];
            end
          else
            begin
              reg546 <= $signed(($unsigned($unsigned(reg520)) ?
                  (-(forvar523 & $signed(wire0))) : $signed((reg505 ^ (reg534 ?
                      reg524 : forvar502)))));
              reg547 <= reg524[(1'h0):(1'h0)];
              reg548 <= {(reg11 <= $unsigned($unsigned($signed(reg496)))),
                  ($signed($signed((8'hae))) < $signed(wire3[(2'h3):(1'h1)]))};
            end
        end
    end
  assign wire551 = $unsigned((~&(~(8'ha9))));
  assign wire552 = forvar491[(3'h4):(2'h3)];
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(reg504)))
        begin
          reg553 = ("S7M0UH5ui" ? (-(~reg14[(4'hb):(3'h7)])) : (~forvar541));
          for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
            begin
              reg555 = $signed((($signed((reg489 ? (8'hbe) : wire1)) ?
                      forvar500 : "agr3") ?
                  ((~&$unsigned(forvar554)) || (~|(8'ha6))) : (reg9[(4'hf):(4'h9)] - (-(!(8'h9f))))));
              reg556 <= (reg6[(5'h12):(4'he)] ~^ reg7[(1'h0):(1'h0)]);
            end
          for (forvar557 = (1'h0); (forvar557 < (3'h4)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 <= (reg546 ? $signed((~$signed(reg529))) : (8'h9e));
              reg559 = (-(($signed((reg542 ? reg504 : reg545)) ?
                      {reg542[(2'h3):(1'h0)], reg525} : (8'hba)) ?
                  ($signed(reg529[(3'h6):(3'h4)]) ?
                      reg492[(4'h8):(3'h5)] : (-forvar514)) : $signed(reg521[(3'h5):(3'h5)])));
              reg560 <= $signed(((8'haa) ?
                  reg511[(4'h9):(3'h5)] : $unsigned($signed(reg520))));
            end
          for (forvar561 = (1'h0); (forvar561 < (1'h0)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 <= reg6[(4'hb):(1'h1)];
              reg563 = ((+$signed(forvar541[(3'h4):(3'h4)])) ?
                  reg560[(5'h10):(4'hf)] : $signed(((reg537[(4'h9):(3'h4)] != $signed(reg501)) ?
                      (^~(reg530 ~^ reg489)) : ($signed(reg507) ?
                          (reg548 & wire552) : (reg550 * reg499)))));
            end
          for (forvar564 = (1'h0); (forvar564 < (3'h4)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 = ({(+reg528[(4'hf):(4'hc)]), forvar491} ?
                  reg559 : (~(($signed((8'ha0)) << $signed(wire552)) ?
                      {""} : (((8'ha1) ? reg563 : (8'hb3)) ~^ (|reg512)))));
              reg566 = $unsigned(reg527[(3'h4):(1'h1)]);
              reg567 = $signed($unsigned(forvar490[(1'h0):(1'h0)]));
              reg568 <= (forvar564[(1'h1):(1'h0)] * (8'had));
              reg569 = forvar541[(2'h2):(1'h1)];
            end
        end
      else
        begin
          for (forvar553 = (1'h0); (forvar553 < (1'h0)); forvar553 = (forvar553 + (1'h1)))
            begin
              reg554 = reg537[(4'hd):(1'h0)];
              reg555 = forvar536[(2'h3):(1'h0)];
              reg556 <= wire60;
              reg557 = forvar490[(2'h2):(1'h1)];
              reg558 = (^~(($signed("IrBYUXoMKzxtPGE2") ?
                      reg535 : (wire551 ?
                          reg9[(4'h8):(2'h3)] : $unsigned(reg543))) ?
                  (reg509[(1'h0):(1'h0)] | forvar491[(2'h2):(2'h2)]) : reg545));
            end
          if ($signed(($unsigned(forvar506) ?
              $unsigned(reg497) : ({(wire2 << reg544),
                  reg520} ^~ {$signed(reg507)}))))
            begin
              reg559 <= $unsigned({{$unsigned(forvar561[(3'h5):(2'h2)]),
                      (~$unsigned((8'ha9)))}});
              reg560 = ($unsigned("w4DXHgsmf59l29") ?
                  (forvar553[(3'h4):(1'h1)] < (reg553[(1'h0):(1'h0)] ?
                      $unsigned({reg567}) : ((^(8'hb1)) && $unsigned(reg503)))) : ((-reg518[(2'h2):(2'h2)]) ?
                      ((!forvar523) ?
                          forvar531[(1'h1):(1'h1)] : (~^$unsigned(reg549))) : (({reg560,
                          reg526} ^~ $signed(forvar516)) <= $unsigned(forvar514))));
              reg561 = (~&wire2[(3'h6):(2'h3)]);
              reg562 <= $signed(($signed($unsigned((reg566 >>> reg510))) ?
                  reg518 : (~|($signed(reg492) <= (reg565 ?
                      forvar561 : reg526)))));
              reg563 <= (forvar554 & (+forvar500));
            end
          else
            begin
              reg559 = ($unsigned({$unsigned((reg567 ?
                      reg495 : reg550))}) && (reg494[(3'h4):(2'h2)] ?
                  "mqduyLtfF3MK" : ($signed({reg568}) ?
                      reg554[(4'hf):(3'h4)] : reg14)));
              reg560 = ({$signed({reg525, (forvar554 ^~ reg558)}),
                      reg539[(4'ha):(4'h8)]} ?
                  reg567[(3'h6):(1'h0)] : {($unsigned(reg537) ?
                          $signed(forvar553[(3'h6):(2'h2)]) : reg532)});
              reg561 = {$unsigned((^~reg499[(1'h1):(1'h0)]))};
              reg562 = {wire487[(3'h4):(2'h2)],
                  ("8iShA0SA" ? $unsigned(reg512) : $unsigned((-reg544)))};
              reg563 = $signed($unsigned(($signed(reg9) >> forvar490)));
            end
          for (forvar564 = (1'h0); (forvar564 < (2'h3)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 = forvar564[(3'h4):(1'h1)];
              reg566 <= ($unsigned(((~^(reg505 ? forvar6 : reg524)) ?
                      forvar500[(4'he):(3'h5)] : $signed((forvar491 <= reg520)))) ?
                  reg550 : reg518);
              reg567 <= (forvar541[(3'h6):(1'h0)] <= $unsigned({(reg557[(3'h4):(2'h3)] ?
                      ((8'hba) + (8'ha5)) : $signed(forvar561))}));
              reg568 = $signed($unsigned((^~($signed(reg547) ?
                  forvar554[(1'h0):(1'h0)] : reg557))));
              reg569 = ($unsigned({((reg518 ~^ forvar517) >= (reg513 ~^ reg569))}) << reg537);
            end
        end
      reg570 <= (^~$unsigned(((8'hb0) ^~ ({reg530} < reg543[(1'h1):(1'h0)]))));
      for (forvar571 = (1'h0); (forvar571 < (2'h3)); forvar571 = (forvar571 + (1'h1)))
        begin
          reg572 <= (((({(8'hab)} ? $signed((8'ha6)) : (forvar541 ~^ (7'h43))) ?
              ($unsigned(wire3) < forvar561[(2'h2):(1'h1)]) : $signed($signed(reg11))) ^ $signed((((8'hbb) | (8'hae)) ?
              {reg550} : (reg13 && (8'ha8))))) | forvar561[(2'h2):(2'h2)]);
          for (forvar573 = (1'h0); (forvar573 < (3'h4)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 <= (((($signed(forvar523) ?
                              $signed(forvar506) : $signed(reg9)) ?
                          ($unsigned(reg534) ?
                              $signed(forvar6) : $signed((8'ha0))) : $unsigned((reg5 ?
                              reg6 : (8'ha0)))) ?
                      reg556 : (8'hb7)) ?
                  reg530 : ((reg549[(1'h1):(1'h1)] ^ reg13) ?
                      (forvar571 << (reg510[(4'ha):(4'ha)] << (~&reg9))) : ($unsigned((-reg499)) && reg539[(5'h10):(3'h6)])));
            end
          if (forvar553)
            begin
              reg575 <= $unsigned("ox");
              reg576 <= $signed(($signed(reg13) ?
                  ((^(forvar506 ?
                      reg495 : reg535)) - {$signed(reg510)}) : reg14[(3'h4):(2'h2)]));
              reg577 <= $unsigned(reg554[(4'hf):(4'hf)]);
              reg578 <= $unsigned((($unsigned({forvar514}) + (~^$signed(wire60))) | (~|(^~(|forvar561)))));
            end
          else
            begin
              reg575 <= forvar514;
              reg576 <= (($unsigned($unsigned((forvar523 ?
                      (8'ha0) : (8'hbb)))) & ($signed((wire0 ?
                      (8'h9c) : (8'hb5))) & reg549)) ?
                  {{((|reg12) == wire4[(1'h0):(1'h0)])},
                      ({forvar573[(4'hc):(3'h7)], (8'hbf)} ?
                          forvar538 : $signed((&reg12)))} : $unsigned(reg534[(4'ha):(3'h4)]));
              reg577 = $signed({reg524[(3'h6):(3'h4)],
                  {(~reg578[(1'h1):(1'h1)])}});
              reg578 = reg558[(1'h0):(1'h0)];
            end
          for (forvar579 = (1'h0); (forvar579 < (3'h4)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 <= "D8QOn1h";
              reg581 <= "GhzQvWPhhu";
              reg582 <= reg492[(4'hf):(4'hd)];
            end
        end
      for (forvar583 = (1'h0); (forvar583 < (1'h0)); forvar583 = (forvar583 + (1'h1)))
        begin
          for (forvar584 = (1'h0); (forvar584 < (3'h4)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 = (reg576 ^~ $signed($signed(((reg532 && reg544) ?
                  forvar502 : $signed(reg537)))));
              reg586 = $signed(($signed(reg549[(2'h2):(1'h0)]) ?
                  $unsigned({{forvar523}}) : (~$unsigned((reg493 ?
                      reg567 : (7'h40))))));
              reg587 = ((+($signed({wire3, (8'hb1)}) ?
                      ({forvar531, reg532} > ((8'hbb) ?
                          (8'hae) : forvar531)) : $signed((~|reg528)))) ?
                  (reg562[(2'h3):(1'h0)] >= $unsigned(((reg544 && wire2) ?
                      reg586 : "kaY"))) : $unsigned(($unsigned({reg501}) >>> $unsigned(forvar523))));
              reg588 <= (^~reg561[(2'h2):(1'h0)]);
            end
          reg589 <= ("F9kNN3" ?
              $signed({{(reg513 <= reg539)}, (~|$signed(reg524))}) : (reg518 ?
                  (8'ha9) : reg586));
          reg590 = {{$unsigned(({reg562} >>> $unsigned((8'hac)))),
                  reg569[(2'h2):(1'h1)]}};
          for (forvar591 = (1'h0); (forvar591 < (1'h0)); forvar591 = (forvar591 + (1'h1)))
            begin
              reg592 <= {reg549[(2'h3):(1'h0)]};
              reg593 <= ($signed((!((reg580 ?
                      wire4 : reg10) | $signed((8'hb2))))) ?
                  reg582[(1'h0):(1'h0)] : $unsigned($unsigned({(~|reg539)})));
              reg594 <= reg587[(4'he):(4'h9)];
            end
          for (forvar595 = (1'h0); (forvar595 < (2'h3)); forvar595 = (forvar595 + (1'h1)))
            begin
              reg596 <= (^~(|reg547));
            end
        end
      for (forvar597 = (1'h0); (forvar597 < (1'h1)); forvar597 = (forvar597 + (1'h1)))
        begin
          for (forvar598 = (1'h0); (forvar598 < (2'h2)); forvar598 = (forvar598 + (1'h1)))
            begin
              reg599 = (~&reg572);
              reg600 <= reg543[(3'h5):(1'h0)];
              reg601 = {(~|{reg494})};
            end
        end
    end
  assign wire602 = (&(~^$unsigned($signed((~reg568)))));
  always
    @(posedge clk) begin
      reg603 <= forvar490;
      reg604 = $unsigned($unsigned({((reg565 > reg596) ?
              (&reg534) : $signed((8'hae)))}));
    end
  module62 modinst606 (.y(wire605), .wire67(reg604), .clk(clk), .wire63(reg501), .wire65(reg548), .wire66(reg562), .wire64(reg545));
  always
    @(posedge clk) begin
      reg607 <= ((&$signed($signed((reg7 >= reg565)))) ?
          {$signed($unsigned((reg554 ? reg495 : forvar573))),
              $unsigned((reg532[(4'hd):(4'ha)] > ((8'hb9) >> reg578)))} : {forvar514});
      for (forvar608 = (1'h0); (forvar608 < (1'h1)); forvar608 = (forvar608 + (1'h1)))
        begin
          reg609 = reg13[(2'h2):(1'h1)];
        end
      for (forvar610 = (1'h0); (forvar610 < (1'h0)); forvar610 = (forvar610 + (1'h1)))
        begin
          for (forvar611 = (1'h0); (forvar611 < (3'h4)); forvar611 = (forvar611 + (1'h1)))
            begin
              reg612 <= $signed(((8'ha2) * (reg511 <= ($unsigned(forvar536) ?
                  (forvar579 ? reg505 : forvar597) : (~^forvar523)))));
              reg613 = reg548[(4'hb):(4'h9)];
            end
          for (forvar614 = (1'h0); (forvar614 < (2'h2)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 = {(reg512 ?
                      {(|$unsigned(reg535)),
                          ((reg586 ? wire552 : reg540) ?
                              (forvar541 - (8'hb5)) : (8'hbb))} : forvar591),
                  $unsigned($unsigned(reg511))};
              reg616 = $unsigned($signed($signed($unsigned((forvar514 && reg522)))));
              reg617 <= reg550[(4'h8):(3'h4)];
            end
          for (forvar618 = (1'h0); (forvar618 < (1'h1)); forvar618 = (forvar618 + (1'h1)))
            begin
              reg619 <= $unsigned({reg580, reg547[(4'hb):(4'hb)]});
              reg620 <= wire2[(2'h3):(2'h2)];
              reg621 <= (($signed(($unsigned(wire605) ?
                      $signed((7'h44)) : $unsigned(reg607))) < (8'hae)) ?
                  {reg535[(3'h7):(3'h6)]} : (reg603 != (($signed(reg515) ?
                      reg603 : reg585) ^~ reg492)));
              reg622 <= reg505;
            end
          for (forvar623 = (1'h0); (forvar623 < (1'h0)); forvar623 = (forvar623 + (1'h1)))
            begin
              reg624 <= ((|($signed((reg620 ? reg581 : reg566)) < ((forvar573 ?
                      forvar538 : reg588) ?
                  (8'ha1) : $unsigned(forvar514)))) + reg562[(4'hf):(3'h4)]);
              reg625 <= ((~&((forvar557[(4'hd):(3'h5)] ?
                      reg582 : $unsigned((7'h41))) == reg498[(2'h3):(1'h0)])) ?
                  (^forvar610) : $unsigned({(reg498 ?
                          reg594[(1'h1):(1'h1)] : {(8'hbf), reg492}),
                      (reg600 ?
                          (reg539 ? reg549 : reg540) : (reg12 ?
                              (8'hb1) : wire552))}));
              reg626 <= (^~$signed(wire602[(1'h1):(1'h0)]));
              reg627 <= (^$signed($signed($signed(forvar618[(4'hd):(4'ha)]))));
              reg628 <= reg14;
            end
          for (forvar629 = (1'h0); (forvar629 < (1'h1)); forvar629 = (forvar629 + (1'h1)))
            begin
              reg630 = reg590[(4'he):(3'h6)];
              reg631 <= $unsigned($unsigned((forvar502 && (wire3[(1'h0):(1'h0)] ?
                  (8'hb8) : {reg580, reg522}))));
            end
        end
    end
  assign wire632 = reg539[(4'hc):(3'h5)];
  always
    @(posedge clk) begin
      if (reg547[(1'h0):(1'h0)])
        begin
          for (forvar633 = (1'h0); (forvar633 < (1'h0)); forvar633 = (forvar633 + (1'h1)))
            begin
              reg634 = ((8'ha6) ? $unsigned($signed((8'hbb))) : "AW");
              reg635 <= reg582;
              reg636 <= reg565[(1'h1):(1'h0)];
            end
          for (forvar637 = (1'h0); (forvar637 < (1'h0)); forvar637 = (forvar637 + (1'h1)))
            begin
              reg638 = reg489;
              reg639 <= $signed({((reg630 ?
                          $signed((8'hb7)) : $unsigned(reg510)) ?
                      $signed(forvar595[(2'h2):(1'h1)]) : $signed((~^(8'hb6))))});
            end
          for (forvar640 = (1'h0); (forvar640 < (3'h4)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 <= (((|$signed("FlXGFw8TLGP9J9")) ?
                      (~|reg529) : forvar573) ?
                  forvar611 : (((+(reg556 ? wire487 : reg601)) ?
                      reg625[(1'h1):(1'h0)] : $unsigned(forvar608)) > $signed($signed(forvar640))));
              reg642 = reg501[(5'h12):(3'h7)];
              reg643 <= "0rvSSF7ysfdayDTg";
              reg644 = $signed((($signed("MQbYYBVk") ?
                  ((reg494 ? (8'hb4) : wire1) ?
                      (~wire605) : {reg642}) : (~^$signed((8'ha8)))) << (~{(+reg492),
                  reg594})));
              reg645 <= {$unsigned((reg580[(2'h2):(2'h2)] <<< {reg578,
                      ((8'hb3) ? reg528 : reg556)})),
                  (forvar502[(1'h0):(1'h0)] ?
                      ((~^(^forvar571)) ?
                          (8'had) : {(reg639 ? forvar553 : reg631),
                              (reg625 ?
                                  forvar618 : reg510)}) : $unsigned("cAKFcMrBDcOTSRg"))};
            end
          for (forvar646 = (1'h0); (forvar646 < (2'h2)); forvar646 = (forvar646 + (1'h1)))
            begin
              reg647 = $unsigned(reg14[(4'hf):(3'h7)]);
              reg648 <= (reg497[(4'h8):(2'h3)] ?
                  (~|$unsigned({$unsigned(reg494),
                      $signed((8'h9f))})) : reg529);
              reg649 <= (reg547[(4'he):(3'h6)] && $unsigned(((-(^reg641)) && $signed((reg565 ?
                  reg533 : reg549)))));
            end
          reg650 = "0CPYw3Xkl67MIaJZk0d";
        end
      else
        begin
          reg633 <= (reg604[(3'h7):(2'h2)] || (($unsigned($signed(forvar629)) >= forvar516[(3'h4):(2'h2)]) || $unsigned(($unsigned(reg532) ~^ (&forvar517)))));
        end
      reg651 = reg649;
      for (forvar652 = (1'h0); (forvar652 < (1'h1)); forvar652 = (forvar652 + (1'h1)))
        begin
          for (forvar653 = (1'h0); (forvar653 < (1'h0)); forvar653 = (forvar653 + (1'h1)))
            begin
              reg654 = $unsigned((reg609[(3'h7):(2'h2)] ?
                  {reg638,
                      ($signed(forvar598) <<< (reg501 ?
                          forvar564 : reg572))} : $unsigned($signed((reg545 >= forvar491)))));
              reg655 = reg604[(4'h9):(3'h5)];
              reg656 <= (reg585 >>> $unsigned(reg599[(3'h5):(2'h2)]));
              reg657 <= $unsigned((reg532 - (8'ha5)));
              reg658 = $signed(forvar491);
            end
          for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = $signed(($signed((forvar611 != reg530[(2'h3):(2'h3)])) & (~reg559)));
            end
          reg661 = reg600[(1'h1):(1'h1)];
        end
      if ("BL3JExsJs77Qlf51P")
        begin
          for (forvar662 = (1'h0); (forvar662 < (2'h2)); forvar662 = (forvar662 + (1'h1)))
            begin
              reg663 <= ({(~$signed(reg6))} ?
                  ({((^forvar571) ? (!forvar541) : (7'h43)),
                          $signed((reg600 == forvar6))} ?
                      (~&{$signed((8'ha0))}) : reg489) : ($signed(reg588[(1'h1):(1'h1)]) || {$unsigned((&reg535)),
                      reg526}));
              reg664 = forvar502;
              reg665 <= reg548[(2'h2):(2'h2)];
              reg666 <= reg587;
            end
          reg667 <= (^$signed($unsigned(reg619)));
          reg668 <= forvar640;
          for (forvar669 = (1'h0); (forvar669 < (2'h2)); forvar669 = (forvar669 + (1'h1)))
            begin
              reg670 <= $signed((({((8'haf) ?
                          (8'had) : (8'hae))} && reg645[(4'h8):(3'h5)]) ?
                  $unsigned({reg664, forvar557}) : (($signed(forvar531) ?
                          $unsigned(reg546) : reg525[(1'h1):(1'h1)]) ?
                      forvar536[(2'h3):(2'h3)] : (!((8'ha0) ?
                          forvar640 : reg520)))));
            end
        end
      else
        begin
          reg662 <= $unsigned((~($signed((~^wire3)) ?
              $unsigned(reg540) : ((-reg542) >> reg532))));
          for (forvar663 = (1'h0); (forvar663 < (2'h3)); forvar663 = (forvar663 + (1'h1)))
            begin
              reg664 <= ($unsigned($unsigned(("y1r05XEGlkJZ3Qg1fIdJ" ?
                      (-reg14) : (forvar591 <= reg600)))) ?
                  (^{(reg498[(2'h2):(1'h1)] < (^reg664))}) : (($unsigned(reg5) ?
                      reg626[(4'he):(4'he)] : {(&reg588),
                          {(8'hb0), (8'hb0)}}) >>> (reg656 ?
                      $unsigned(reg616) : ($signed(reg616) ?
                          reg645 : {reg624, reg545}))));
            end
          for (forvar665 = (1'h0); (forvar665 < (1'h1)); forvar665 = (forvar665 + (1'h1)))
            begin
              reg666 = $unsigned(reg501[(1'h0):(1'h0)]);
              reg667 <= $signed((~^(wire632 ?
                  ((^reg512) <<< (reg496 ?
                      reg537 : (8'hb6))) : forvar6[(4'h9):(2'h2)])));
            end
        end
    end
  assign wire671 = forvar623;
  module62 modinst673 (wire672, clk, reg535, forvar637, reg522, forvar561, forvar608);
  always
    @(posedge clk) begin
      for (forvar674 = (1'h0); (forvar674 < (2'h3)); forvar674 = (forvar674 + (1'h1)))
        begin
          reg675 = ({wire2, (^~$signed((reg613 != reg661)))} ?
              $signed(reg616[(3'h4):(2'h3)]) : reg582[(2'h3):(2'h3)]);
        end
    end
  assign wire676 = reg570;
  module324 modinst678 (wire677, clk, reg675, reg627, reg633, reg526);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module62  (y, clk, wire63, wire64, wire65, wire66, wire67);
  output wire [(32'h594):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire63;
  input wire signed [(4'hd):(1'h0)] wire64;
  input wire signed [(4'he):(1'h0)] wire65;
  input wire signed [(5'h15):(1'h0)] wire66;
  input wire signed [(4'hc):(1'h0)] wire67;
  reg [(3'h5):(1'h0)] reg485 = (1'h0);
  reg [(4'he):(1'h0)] forvar480 = (1'h0);
  reg signed [(4'he):(1'h0)] reg486 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar485 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg483 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg482 = (1'h0);
  reg [(3'h6):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg480 = (1'h0);
  reg [(3'h6):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar477 = (1'h0);
  reg [(5'h10):(1'h0)] reg476 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar475 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar474 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg473 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg471 = (1'h0);
  reg [(4'hb):(1'h0)] reg470 = (1'h0);
  reg [(3'h5):(1'h0)] reg469 = (1'h0);
  reg [(4'hb):(1'h0)] forvar468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg467 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg466 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg465 = (1'h0);
  reg [(4'h9):(1'h0)] reg464 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg463 = (1'h0);
  reg [(4'h8):(1'h0)] reg462 = (1'h0);
  reg [(3'h5):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg460 = (1'h0);
  reg [(4'ha):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar458 = (1'h0);
  reg [(4'h8):(1'h0)] forvar457 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg456 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire453;
  wire [(4'hc):(1'h0)] wire323;
  reg signed [(5'h11):(1'h0)] reg322 = (1'h0);
  reg [(5'h14):(1'h0)] forvar321 = (1'h0);
  reg [(3'h7):(1'h0)] forvar320 = (1'h0);
  reg [(3'h4):(1'h0)] reg319 = (1'h0);
  reg [(3'h7):(1'h0)] reg318 = (1'h0);
  reg [(3'h5):(1'h0)] reg317 = (1'h0);
  reg [(5'h14):(1'h0)] reg316 = (1'h0);
  reg [(4'h9):(1'h0)] reg315 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar314 = (1'h0);
  reg [(4'hb):(1'h0)] reg313 = (1'h0);
  reg [(4'hc):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg310 = (1'h0);
  reg [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar306 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg305 = (1'h0);
  reg [(3'h5):(1'h0)] reg304 = (1'h0);
  reg [(4'he):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg300 = (1'h0);
  reg [(5'h11):(1'h0)] forvar299 = (1'h0);
  reg [(2'h3):(1'h0)] reg298 = (1'h0);
  wire [(3'h4):(1'h0)] wire297;
  wire signed [(2'h2):(1'h0)] wire296;
  reg signed [(3'h5):(1'h0)] reg295 = (1'h0);
  reg [(4'he):(1'h0)] reg294 = (1'h0);
  reg [(5'h13):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg290 = (1'h0);
  reg [(2'h2):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg287 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg286 = (1'h0);
  reg [(4'he):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar284 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg283 = (1'h0);
  reg signed [(4'he):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg281 = (1'h0);
  reg [(4'hc):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg279 = (1'h0);
  reg [(3'h7):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg277 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar276 = (1'h0);
  reg signed [(4'he):(1'h0)] reg275 = (1'h0);
  reg [(5'h10):(1'h0)] reg274 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg273 = (1'h0);
  reg [(3'h6):(1'h0)] reg272 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar271 = (1'h0);
  reg signed [(4'he):(1'h0)] reg270 = (1'h0);
  reg [(5'h14):(1'h0)] forvar269 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg266 = (1'h0);
  reg [(5'h10):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg264 = (1'h0);
  reg [(4'hb):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] reg262 = (1'h0);
  reg [(4'hf):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar260 = (1'h0);
  reg [(5'h11):(1'h0)] forvar251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg250 = (1'h0);
  reg signed [(4'he):(1'h0)] reg259 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg258 = (1'h0);
  reg [(4'hf):(1'h0)] reg257 = (1'h0);
  reg [(4'hb):(1'h0)] forvar256 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg254 = (1'h0);
  reg [(4'he):(1'h0)] reg253 = (1'h0);
  reg [(5'h15):(1'h0)] reg252 = (1'h0);
  reg [(4'h8):(1'h0)] reg251 = (1'h0);
  reg [(3'h7):(1'h0)] forvar250 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg248 = (1'h0);
  reg [(5'h15):(1'h0)] reg247 = (1'h0);
  reg [(5'h13):(1'h0)] reg246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg245 = (1'h0);
  reg [(3'h7):(1'h0)] reg244 = (1'h0);
  reg [(5'h15):(1'h0)] forvar243 = (1'h0);
  reg [(4'hf):(1'h0)] reg242 = (1'h0);
  reg [(5'h12):(1'h0)] reg241 = (1'h0);
  wire [(3'h5):(1'h0)] wire240;
  wire signed [(5'h14):(1'h0)] wire68;
  wire [(4'h9):(1'h0)] wire69;
  wire signed [(5'h14):(1'h0)] wire70;
  wire signed [(4'ha):(1'h0)] wire238;
  assign y = {reg485,
                 forvar480,
                 reg486,
                 forvar485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 forvar477,
                 reg476,
                 forvar475,
                 forvar474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 forvar468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 forvar458,
                 forvar457,
                 reg456,
                 reg455,
                 wire453,
                 wire323,
                 reg322,
                 forvar321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 forvar314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 forvar306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 forvar299,
                 reg298,
                 wire297,
                 wire296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 forvar276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 forvar271,
                 reg270,
                 forvar269,
                 reg268,
                 forvar267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 forvar260,
                 forvar251,
                 reg250,
                 reg259,
                 reg258,
                 reg257,
                 forvar256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 forvar250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 forvar243,
                 reg242,
                 reg241,
                 wire240,
                 wire68,
                 wire69,
                 wire70,
                 wire238,
                 (1'h0)};
  assign wire68 = ($unsigned($unsigned(($unsigned(wire65) >> (~|wire67)))) && ($unsigned({{wire63}}) >= $unsigned($unsigned($signed(wire67)))));
  assign wire69 = (("0ElCIHih8wX" ?
                      wire63 : ($signed(((8'hbc) + (8'hb5))) ^~ ({wire66} * wire64[(3'h6):(3'h5)]))) >>> (((wire64[(3'h4):(1'h0)] ?
                          (&wire65) : $unsigned(wire66)) ?
                      wire64 : ((wire68 ~^ wire65) ^~ (wire67 & wire67))) << $signed($signed(wire64))));
  assign wire70 = (~|wire69[(2'h2):(1'h0)]);
  module71 modinst239 (wire238, clk, wire68, wire63, wire66, wire67, wire64);
  assign wire240 = wire63;
  always
    @(posedge clk) begin
      reg241 = $signed(wire240);
      reg242 <= wire67;
      for (forvar243 = (1'h0); (forvar243 < (1'h1)); forvar243 = (forvar243 + (1'h1)))
        begin
          if (wire66)
            begin
              reg244 <= (((($signed(wire69) ~^ reg242[(3'h5):(3'h4)]) ?
                          ((wire238 <<< wire63) ?
                              wire240[(3'h4):(2'h3)] : (8'hb3)) : $signed(wire240[(2'h2):(1'h0)])) ?
                      forvar243 : wire65) ?
                  $unsigned((((reg241 <<< wire63) & $signed((8'hb4))) & reg242[(4'h8):(2'h2)])) : wire63);
              reg245 = wire67;
              reg246 = ($signed($unsigned((wire238 - wire240[(1'h1):(1'h0)]))) ?
                  (((&(&wire66)) ?
                      $unsigned((wire66 ~^ wire67)) : (wire67 + $signed(reg242))) <= (~&("6Bdd7IlSzAkGGSH" | "pHB"))) : $unsigned(wire67[(3'h7):(3'h5)]));
              reg247 = reg244;
            end
          else
            begin
              reg244 = wire66;
            end
          reg248 = (-("J4ZAHZmlhdhU7" ?
              (8'ha4) : $signed(((wire63 ? wire238 : forvar243) ?
                  reg244 : (^wire66)))));
        end
      reg249 = {wire69[(3'h5):(3'h5)],
          ((($unsigned((8'ha1)) ?
              (wire68 ? forvar243 : reg246) : (reg244 ?
                  wire70 : reg241)) < $signed(((8'ha1) ?
              (8'hac) : (8'hb5)))) ~^ (wire63[(3'h4):(1'h1)] && reg242))};
      if ("d0o")
        begin
          for (forvar250 = (1'h0); (forvar250 < (1'h0)); forvar250 = (forvar250 + (1'h1)))
            begin
              reg251 <= $signed({(&(reg244[(2'h3):(2'h3)] ?
                      $unsigned((8'hb1)) : "0")),
                  ({(reg249 ?
                          reg244 : forvar250)} || $unsigned((wire65 <= reg245)))});
              reg252 <= (!$signed((!{((8'hb6) ? reg246 : wire64)})));
              reg253 = ("0qH51GM" ?
                  $signed({((reg249 == wire67) >= {reg242, reg252}),
                      $signed(wire69)}) : $unsigned((wire66[(5'h12):(4'he)] ?
                      $unsigned((wire68 ?
                          wire65 : wire240)) : {wire63[(4'hc):(3'h6)]})));
              reg254 = wire240[(3'h4):(1'h1)];
              reg255 <= (((-$signed(reg254[(4'h8):(1'h0)])) && (wire66[(4'hc):(2'h2)] ?
                  $signed({(8'hae)}) : wire64)) || $unsigned($unsigned((+(!reg248)))));
            end
          for (forvar256 = (1'h0); (forvar256 < (1'h1)); forvar256 = (forvar256 + (1'h1)))
            begin
              reg257 <= $unsigned($unsigned(wire240));
              reg258 = (~^wire67);
              reg259 <= $unsigned(wire70);
            end
        end
      else
        begin
          reg250 <= (!reg255[(2'h2):(1'h0)]);
          for (forvar251 = (1'h0); (forvar251 < (2'h3)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 <= $unsigned((7'h41));
              reg253 <= wire68[(5'h12):(3'h6)];
              reg254 <= wire65;
              reg255 <= $signed(($signed({((8'h9e) ? reg250 : (8'hb5)),
                  $unsigned((8'hb2))}) < forvar243));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar260 = (1'h0); (forvar260 < (1'h1)); forvar260 = (forvar260 + (1'h1)))
        begin
          if ((reg247[(2'h2):(1'h0)] ?
              $signed(reg251[(1'h0):(1'h0)]) : $unsigned((~^(reg241[(4'ha):(4'h9)] + $signed(forvar256))))))
            begin
              reg261 <= ($signed({wire69[(3'h6):(1'h0)],
                  $signed({wire64})}) >= reg246[(5'h10):(4'hd)]);
              reg262 <= "eEfv";
              reg263 <= (((8'hbf) ?
                      reg250 : (^(((8'hb3) >>> reg262) << (&wire65)))) ?
                  wire64[(3'h6):(3'h4)] : ((reg254[(3'h5):(2'h3)] <<< (8'hb8)) ^ (&(8'ha9))));
            end
          else
            begin
              reg261 = ({$unsigned(reg258)} ?
                  reg259 : (~&({wire240[(2'h2):(1'h0)],
                      (wire65 ? wire240 : wire65)} == (~$signed(forvar251)))));
              reg262 <= $unsigned((!((8'hb8) | ((forvar250 ? reg255 : (8'haf)) ?
                  (~|reg248) : {reg245, reg263}))));
              reg263 <= $signed(wire64);
              reg264 <= ((+(8'hbf)) ?
                  $signed($unsigned({{wire240, wire238},
                      $unsigned(reg255)})) : wire63[(4'hc):(3'h5)]);
            end
          reg265 <= (&reg252);
        end
      reg266 = $unsigned(reg261[(1'h1):(1'h0)]);
      for (forvar267 = (1'h0); (forvar267 < (1'h0)); forvar267 = (forvar267 + (1'h1)))
        begin
          reg268 <= reg262[(2'h2):(1'h0)];
          for (forvar269 = (1'h0); (forvar269 < (3'h4)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 <= $signed({$unsigned($signed((reg263 & wire240))),
                  ((reg250 + {(8'hab),
                      (8'hb6)}) != (forvar243[(1'h1):(1'h0)] ^~ $signed(forvar267)))});
            end
          for (forvar271 = (1'h0); (forvar271 < (2'h2)); forvar271 = (forvar271 + (1'h1)))
            begin
              reg272 <= "Y5o2x0";
              reg273 = {reg264[(4'hb):(3'h7)], forvar243};
              reg274 <= (^~{($unsigned(reg244[(1'h0):(1'h0)]) << reg252[(4'hf):(1'h0)])});
              reg275 <= {$signed((~^({reg255, wire70} ?
                      (reg254 ^~ reg242) : (forvar267 || wire66)))),
                  $unsigned((-{((8'hb5) ? reg253 : (7'h43))}))};
            end
          for (forvar276 = (1'h0); (forvar276 < (1'h1)); forvar276 = (forvar276 + (1'h1)))
            begin
              reg277 <= reg250;
              reg278 = $unsigned((((+(wire68 ? (8'h9f) : reg266)) ?
                      "TZ1EXfC5eDvZ0q" : ((^~reg277) ?
                          (reg265 == wire240) : wire67)) ?
                  $signed((~&(reg262 < (7'h41)))) : $signed((~wire66[(4'ha):(1'h0)]))));
              reg279 = (|(~((!reg250) ?
                  forvar269[(2'h3):(2'h2)] : reg255[(2'h2):(1'h0)])));
            end
          if (((^~reg265[(4'h9):(1'h0)]) << wire69))
            begin
              reg280 <= $signed(reg273);
              reg281 = ($unsigned(wire64[(1'h1):(1'h0)]) ?
                  {((^{reg265, reg257}) ? (8'ha8) : wire70[(5'h12):(5'h12)]),
                      $unsigned((((8'hb6) + reg266) ?
                          (wire238 * reg273) : (reg251 + reg252)))} : ({$signed((reg248 * wire238))} ?
                      {(!(!(8'hb1))),
                          $unsigned(((7'h41) * wire238))} : reg263[(4'ha):(3'h6)]));
              reg282 <= $unsigned(forvar269);
            end
          else
            begin
              reg280 <= (((forvar256 & wire238) - (((^~wire64) ?
                          (reg263 || wire66) : (reg254 ^ reg258)) ?
                      reg272[(2'h3):(2'h2)] : $signed((reg247 ^~ reg275)))) ?
                  (reg252[(4'hd):(1'h1)] ?
                      wire65[(1'h1):(1'h0)] : $signed((~|wire63))) : $unsigned($unsigned(forvar250[(1'h0):(1'h0)])));
              reg281 <= ({reg261} ?
                  $signed(forvar276) : $unsigned((~($signed(reg246) ?
                      $unsigned(reg242) : $unsigned((7'h43))))));
              reg282 <= reg265;
              reg283 = ((7'h40) == $signed($signed((reg241[(3'h6):(1'h0)] ^~ $signed(forvar251)))));
            end
        end
      for (forvar284 = (1'h0); (forvar284 < (1'h0)); forvar284 = (forvar284 + (1'h1)))
        begin
          reg285 <= $unsigned("Uq6");
          if ($signed($unsigned(($unsigned(((7'h42) * forvar276)) >> {reg242,
              (reg251 ? wire69 : forvar276)}))))
            begin
              reg286 <= reg265[(4'h9):(4'h8)];
              reg287 <= reg272[(2'h2):(1'h1)];
              reg288 <= $unsigned($unsigned((wire64 ?
                  {wire68[(5'h11):(3'h5)],
                      "dT9ReiKbSJO"} : reg244[(1'h1):(1'h1)])));
              reg289 <= (~&reg274[(4'hb):(4'h8)]);
            end
          else
            begin
              reg286 <= (reg263[(2'h2):(2'h2)] ?
                  $signed($signed("4QphFcy")) : ((($signed(reg266) ?
                          {reg255} : reg270) ^ ($signed(reg241) ^~ ((8'hae) > reg258))) ?
                      {$unsigned($unsigned((8'hb2))),
                          (8'ha0)} : reg273[(1'h1):(1'h1)]));
            end
          reg290 <= $signed(forvar284);
          if ((|reg279[(5'h13):(3'h4)]))
            begin
              reg291 <= ((+$signed($signed((^forvar250)))) ?
                  (^~((+$unsigned(forvar284)) & ((~reg263) && $unsigned(reg262)))) : $unsigned(wire238));
              reg292 = (reg249[(2'h3):(2'h3)] <= (($signed({forvar250,
                          reg282}) ?
                      (reg266[(3'h7):(2'h3)] ?
                          reg265 : forvar250) : ("m50afalf4OEDZp" ?
                          (wire68 ? forvar250 : reg242) : $unsigned(reg285))) ?
                  ($unsigned(reg242[(2'h3):(1'h1)]) ?
                      (reg251 << (forvar267 == reg275)) : (~|forvar284[(3'h5):(2'h3)])) : $signed($unsigned(((8'ha7) * reg290)))));
              reg293 <= ($signed(((8'hba) - $signed(reg289))) ^~ $signed(($unsigned(reg266[(3'h6):(1'h0)]) <<< wire240)));
              reg294 <= reg258;
              reg295 <= {((|((&reg275) << reg290)) ?
                      (&"CnHRYTPM") : ($unsigned((wire240 ? (7'h40) : reg293)) ?
                          ((reg279 ? reg279 : reg259) ?
                              (reg291 <<< reg273) : ((8'hb8) ?
                                  reg288 : forvar267)) : ((reg242 - reg288) ?
                              (reg257 ^ reg277) : $unsigned(wire64))))};
            end
          else
            begin
              reg291 <= (~&"gIBMOGOq8csiiOqfy6Sf");
              reg292 = $signed(forvar260);
            end
        end
    end
  assign wire296 = reg259;
  assign wire297 = {({$unsigned((forvar271 ? reg272 : reg259)),
                               reg261[(3'h4):(1'h1)]} ?
                           ($unsigned({reg255}) <= $unsigned(((8'hb3) << reg244))) : ((8'ha0) ?
                               $unsigned($unsigned(reg244)) : reg253[(3'h5):(2'h3)])),
                       (($unsigned((forvar256 << (8'ha0))) >= $unsigned($signed(wire68))) ~^ (-(reg244 ?
                           wire70[(5'h14):(4'ha)] : (&(7'h42)))))};
  always
    @(posedge clk) begin
      reg298 = "t";
      for (forvar299 = (1'h0); (forvar299 < (1'h1)); forvar299 = (forvar299 + (1'h1)))
        begin
          if (($unsigned(reg282[(2'h3):(2'h3)]) && ((~^((reg263 + reg287) ?
                  ((8'hba) ? wire297 : forvar267) : "YXFmpi")) ?
              (^~wire67) : {{((8'hbd) && reg295), forvar243[(1'h0):(1'h0)]},
                  ((wire68 << reg265) ?
                      (forvar267 ? reg293 : reg291) : (&reg248))})))
            begin
              reg300 = (-$unsigned($unsigned($signed($signed(reg278)))));
            end
          else
            begin
              reg300 <= (reg291 >>> {(reg281[(3'h4):(3'h4)] ?
                      (reg254 == wire66[(5'h11):(3'h6)]) : (+$signed(wire66)))});
              reg301 = wire297;
              reg302 <= $unsigned($unsigned($unsigned(({reg254,
                  reg282} > reg278[(1'h0):(1'h0)]))));
              reg303 <= ((reg293[(4'hc):(3'h6)] & $signed($signed($signed((8'h9d))))) == (&wire297[(1'h0):(1'h0)]));
              reg304 = ("ry4tla3XGyHWyK" ? (+(^~(^{wire70}))) : reg298);
            end
        end
      reg305 = (forvar250[(3'h5):(3'h5)] ?
          {(((reg292 == reg259) ?
                  $unsigned(reg250) : {reg278}) != reg252[(4'h8):(3'h4)])} : (&$unsigned(reg291[(5'h13):(5'h10)])));
      for (forvar306 = (1'h0); (forvar306 < (2'h3)); forvar306 = (forvar306 + (1'h1)))
        begin
          if (wire64)
            begin
              reg307 = reg294[(4'h8):(3'h4)];
              reg308 <= reg272;
              reg309 <= ($unsigned((reg244 << ($unsigned(reg257) ?
                  ((8'hb3) + forvar267) : reg248[(1'h0):(1'h0)]))) & {reg287[(3'h6):(3'h4)]});
            end
          else
            begin
              reg307 = reg304;
              reg308 = {$signed((^~(reg250[(2'h2):(1'h1)] ?
                      $unsigned(reg259) : $unsigned(reg303)))),
                  (reg274 >>> {{(~|reg257)}})};
              reg309 <= (~&(|(wire68 == reg287[(3'h6):(3'h5)])));
            end
          reg310 <= (reg288 || reg253);
        end
    end
  always
    @(posedge clk) begin
      reg311 = $signed((($unsigned(reg295[(3'h5):(2'h2)]) << forvar306) != (8'ha4)));
      reg312 <= ("K" || $signed(("VF7rce2wiifX7N" ?
          $signed($signed(reg311)) : "48R")));
      reg313 <= (!({{$unsigned((8'hb6)), $unsigned(reg274)}, reg279} ?
          $unsigned(($signed(reg281) + $unsigned(wire297))) : $unsigned("cIp8ThVZ")));
      if ($signed((!$signed(forvar267))))
        begin
          for (forvar314 = (1'h0); (forvar314 < (2'h3)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg315 <= (!((^~forvar243) ?
                  (reg304[(1'h1):(1'h1)] ?
                      $unsigned($signed(reg278)) : ({(8'hb3), forvar276} ?
                          reg282 : "")) : (reg268[(1'h0):(1'h0)] != ($signed(reg278) || $signed(reg247)))));
              reg316 <= ($unsigned("21u") ^ $unsigned((&$unsigned(reg298[(2'h3):(2'h2)]))));
              reg317 <= $signed($signed(($signed((!reg253)) >= forvar256[(1'h1):(1'h0)])));
              reg318 = ((reg304 ?
                      reg281[(2'h2):(1'h0)] : $unsigned(((-reg265) ?
                          reg316[(4'hd):(4'h8)] : (^(8'h9f))))) ?
                  wire64 : (~{$signed(wire66[(1'h0):(1'h0)]),
                      ((-wire240) ?
                          (reg283 <<< forvar299) : (reg289 >= reg252))}));
              reg319 <= ($signed(((reg290 ? (&(8'ha5)) : {reg308, reg263}) ?
                  $unsigned($signed(forvar276)) : "k")) + $unsigned((reg317 + ((wire296 ?
                      (8'ha7) : forvar256) ?
                  (reg274 ? reg242 : reg303) : (reg274 & (8'h9f))))));
            end
        end
      else
        begin
          for (forvar314 = (1'h0); (forvar314 < (3'h4)); forvar314 = (forvar314 + (1'h1)))
            begin
              reg315 <= ((+(&(reg308 ?
                      (^forvar243) : (reg248 ? (8'hbe) : reg247)))) ?
                  {$signed(reg288),
                      ($unsigned((~&reg263)) ?
                          $signed(reg288) : ((wire66 ?
                              reg317 : reg275) != $signed(reg305)))} : reg253[(2'h2):(2'h2)]);
            end
          reg316 = ({$signed((^forvar306))} << (reg257[(3'h7):(3'h4)] != ((+reg248) ?
              reg246 : {$unsigned((8'ha7))})));
        end
      for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
        begin
          for (forvar321 = (1'h0); (forvar321 < (1'h1)); forvar321 = (forvar321 + (1'h1)))
            begin
              reg322 <= forvar299[(3'h7):(1'h0)];
            end
        end
    end
  assign wire323 = {$signed({$unsigned(((7'h40) > reg242)),
                           ((reg322 != reg312) ^~ $unsigned(reg293))})};
  module324 modinst454 (.wire326(reg280), .y(wire453), .clk(clk), .wire325(reg318), .wire327(reg270), .wire328(reg245));
  always
    @(posedge clk) begin
      reg455 = $signed((8'ha7));
      reg456 <= (wire63 ?
          (~|$unsigned((((8'ha8) ? reg291 : wire67) ?
              reg293[(4'ha):(2'h2)] : {reg315}))) : $unsigned(reg290[(4'he):(3'h6)]));
      for (forvar457 = (1'h0); (forvar457 < (3'h4)); forvar457 = (forvar457 + (1'h1)))
        begin
          for (forvar458 = (1'h0); (forvar458 < (2'h2)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 = forvar276[(3'h5):(3'h4)];
              reg460 = {(^$signed(reg241))};
              reg461 <= forvar243[(3'h4):(3'h4)];
              reg462 <= reg279[(1'h1):(1'h1)];
            end
          if ((reg318 ?
              (|reg286) : (((reg310[(1'h1):(1'h1)] ?
                      reg241[(5'h10):(3'h5)] : {reg300, forvar251}) ?
                  ($signed(forvar284) ?
                      wire297[(2'h3):(1'h1)] : (reg319 ?
                          reg460 : reg281)) : (((8'ha0) ? (8'hab) : reg280) ?
                      (reg303 < reg272) : {reg298})) > (forvar458 * (8'hbf)))))
            begin
              reg463 <= $unsigned(reg273[(2'h2):(1'h0)]);
              reg464 <= reg265;
              reg465 <= reg255;
              reg466 <= (|(7'h41));
              reg467 <= reg266;
            end
          else
            begin
              reg463 <= (^~reg307[(1'h0):(1'h0)]);
              reg464 <= $signed((~(8'ha2)));
              reg465 <= ((reg250 == {((-reg317) > $unsigned(wire63))}) ~^ ({$unsigned((~reg465)),
                      (-(^reg254))} ?
                  reg262 : $unsigned((~|(^reg254)))));
              reg466 = (8'ha3);
              reg467 <= {((^~$unsigned((reg322 >= reg459))) ?
                      $signed((~(8'ha6))) : (~&(((8'hae) ?
                          reg455 : reg312) > $unsigned(reg272)))),
                  $unsigned((^forvar251[(4'ha):(2'h3)]))};
            end
          for (forvar468 = (1'h0); (forvar468 < (2'h3)); forvar468 = (forvar468 + (1'h1)))
            begin
              reg469 = reg313;
              reg470 <= ((reg466[(3'h7):(2'h2)] ?
                  {$unsigned(reg272),
                      wire64[(1'h0):(1'h0)]} : "DKly0") | $unsigned($unsigned((^$signed(reg245)))));
              reg471 <= (($signed((|$signed(reg247))) ?
                  (wire297[(1'h0):(1'h0)] ?
                      $signed(reg273[(1'h1):(1'h0)]) : (~^reg266[(1'h1):(1'h1)])) : $unsigned(($signed(reg273) ?
                      (^~reg281) : (~^wire65)))) << $signed($signed((&$signed(reg302)))));
              reg472 <= reg291;
            end
          reg473 = (|$signed((reg270 + forvar314[(4'h8):(3'h5)])));
        end
      for (forvar474 = (1'h0); (forvar474 < (1'h1)); forvar474 = (forvar474 + (1'h1)))
        begin
          for (forvar475 = (1'h0); (forvar475 < (3'h4)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 <= $signed(reg463);
            end
          for (forvar477 = (1'h0); (forvar477 < (3'h4)); forvar477 = (forvar477 + (1'h1)))
            begin
              reg478 <= wire297;
              reg479 <= ((forvar256[(3'h6):(2'h2)] == (reg281 ?
                  forvar256 : (~|(forvar267 * reg281)))) >>> reg250[(2'h3):(2'h3)]);
            end
        end
      if ($unsigned({$signed(reg251[(3'h5):(3'h4)])}))
        begin
          if (reg247[(1'h1):(1'h1)])
            begin
              reg480 = {reg308,
                  ((reg286 ?
                          reg272 : ((!reg248) ?
                              {reg301} : (wire240 ? wire65 : reg255))) ?
                      (^~forvar475) : $signed((reg264 ?
                          ((8'ha7) >> reg469) : (reg244 > reg272))))};
              reg481 <= $unsigned((8'ha4));
              reg482 <= ($unsigned(((!$unsigned(reg264)) <<< $unsigned($signed(reg308)))) <= reg310[(1'h0):(1'h0)]);
            end
          else
            begin
              reg480 <= $signed(($unsigned((~^((8'ha9) ?
                  reg293 : reg460))) ~^ forvar468[(4'hb):(1'h1)]));
              reg481 <= {((($unsigned(forvar243) ?
                      ((8'ha3) ?
                          reg293 : forvar251) : (!reg287)) >>> reg270[(4'he):(1'h1)]) <= wire297)};
              reg482 <= reg466[(1'h0):(1'h0)];
              reg483 = reg290[(4'hf):(4'he)];
              reg484 <= (~|$signed({reg322[(4'hf):(2'h3)], reg294}));
            end
          for (forvar485 = (1'h0); (forvar485 < (3'h4)); forvar485 = (forvar485 + (1'h1)))
            begin
              reg486 <= $unsigned((wire238[(4'h8):(2'h2)] ?
                  forvar260 : $signed($unsigned(reg287[(3'h7):(1'h1)]))));
            end
        end
      else
        begin
          for (forvar480 = (1'h0); (forvar480 < (2'h2)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 = forvar243[(4'ha):(4'ha)];
              reg482 <= reg277;
              reg483 <= (((forvar468[(4'h8):(2'h2)] ?
                      ((|reg246) ?
                          $unsigned(reg301) : $unsigned(reg483)) : $unsigned($signed(reg258))) == ((+(^~(8'had))) ?
                      $signed({reg300}) : (wire68[(4'hb):(2'h2)] ?
                          (~|reg253) : forvar458))) ?
                  (~|(reg258 ?
                      $unsigned((~|reg255)) : ($signed(reg315) ?
                          (^reg286) : (forvar475 < (8'hb7))))) : ((wire64[(4'h8):(2'h2)] >>> $unsigned(reg247[(4'h9):(2'h2)])) ?
                      "99DQqUYqPvNoX" : $signed($signed(reg285))));
              reg484 <= reg290[(4'h8):(1'h1)];
            end
          reg485 <= forvar243[(5'h14):(4'h8)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module15
#( parameter param58 = {{(~(((8'h9e) ? (8'ha0) : (8'hbd)) ? ((8'h9f) ^ (8'ha9)) : ((8'hb8) & (7'h44))))}}
, parameter param59 = {param58, ((((param58 ? param58 : param58) << {(8'hbf)}) <= param58) ? param58 : param58)} )
(y, clk, wire20, wire19, wire18, wire17, wire16);
  output wire [(32'h1da):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire20;
  input wire [(4'ha):(1'h0)] wire19;
  input wire [(5'h10):(1'h0)] wire18;
  input wire signed [(5'h13):(1'h0)] wire17;
  input wire signed [(2'h2):(1'h0)] wire16;
  wire signed [(4'hc):(1'h0)] wire57;
  wire [(5'h13):(1'h0)] wire56;
  reg [(5'h11):(1'h0)] reg55 = (1'h0);
  reg [(2'h3):(1'h0)] forvar54 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar53 = (1'h0);
  reg [(5'h13):(1'h0)] reg52 = (1'h0);
  reg [(3'h7):(1'h0)] reg51 = (1'h0);
  reg [(3'h5):(1'h0)] reg50 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar48 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar47 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar42 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg38 = (1'h0);
  reg [(5'h13):(1'h0)] forvar35 = (1'h0);
  reg [(5'h10):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg44 = (1'h0);
  reg [(2'h3):(1'h0)] reg43 = (1'h0);
  reg [(2'h3):(1'h0)] reg42 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg41 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar38 = (1'h0);
  reg [(2'h3):(1'h0)] reg37 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg35 = (1'h0);
  reg [(5'h14):(1'h0)] reg34 = (1'h0);
  reg [(5'h15):(1'h0)] reg33 = (1'h0);
  reg [(3'h4):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg30 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar29 = (1'h0);
  reg [(2'h2):(1'h0)] reg28 = (1'h0);
  reg [(3'h6):(1'h0)] forvar27 = (1'h0);
  reg [(3'h7):(1'h0)] reg26 = (1'h0);
  reg [(5'h12):(1'h0)] forvar25 = (1'h0);
  reg [(5'h14):(1'h0)] reg24 = (1'h0);
  reg [(2'h2):(1'h0)] reg23 = (1'h0);
  wire [(5'h15):(1'h0)] wire22;
  wire [(5'h13):(1'h0)] wire21;
  assign y = {wire57,
                 wire56,
                 reg55,
                 forvar54,
                 forvar53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 forvar48,
                 forvar47,
                 forvar42,
                 reg38,
                 forvar35,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 forvar38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 reg28,
                 forvar27,
                 reg26,
                 forvar25,
                 reg24,
                 reg23,
                 wire22,
                 wire21,
                 (1'h0)};
  assign wire21 = wire16;
  assign wire22 = wire18;
  always
    @(posedge clk) begin
      reg23 = wire17;
      reg24 = $signed($unsigned({((^wire21) <<< (^~(8'haa)))}));
      for (forvar25 = (1'h0); (forvar25 < (1'h1)); forvar25 = (forvar25 + (1'h1)))
        begin
          reg26 <= $signed((($unsigned(reg23[(1'h1):(1'h0)]) ?
                  "" : wire20[(3'h7):(3'h7)]) ?
              ((((8'hbb) ? wire20 : wire22) ?
                      (wire16 != reg24) : {wire22, wire18}) ?
                  ("c3aZobCBl8b1XylvSpZ" != wire20) : (((8'ha6) ?
                          reg24 : (8'hbf)) ?
                      wire21[(4'hf):(4'hf)] : (wire17 ?
                          wire17 : wire16))) : ("zwPdZb09oXwQ" ?
                  (~|(8'hb6)) : ((|(8'hb6)) + (|wire16)))));
          for (forvar27 = (1'h0); (forvar27 < (1'h0)); forvar27 = (forvar27 + (1'h1)))
            begin
              reg28 <= (~&($unsigned(wire22) >= reg23[(1'h0):(1'h0)]));
            end
          for (forvar29 = (1'h0); (forvar29 < (2'h2)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 = wire19[(3'h4):(3'h4)];
              reg31 <= $unsigned((($signed((8'ha7)) ?
                  reg26 : {{reg26, wire20}}) >> ((!$signed(forvar27)) ?
                  reg30[(1'h0):(1'h0)] : (|"h8xVJZ3Xz815s1RSPnok"))));
            end
        end
      reg32 <= ({$unsigned($signed(((7'h43) ? wire21 : (8'h9d)))),
          wire17[(3'h5):(1'h1)]} & reg24);
    end
  always
    @(posedge clk) begin
      reg33 = wire20;
      if ((7'h40))
        begin
          if ((~|reg30))
            begin
              reg34 <= (|$unsigned(({$unsigned(reg23), $signed(reg28)} ?
                  ((8'ha9) ?
                      $signed(wire22) : wire21[(5'h13):(5'h13)]) : $unsigned($unsigned((8'hb4))))));
              reg35 <= (7'h40);
            end
          else
            begin
              reg34 <= (wire16[(1'h1):(1'h1)] >>> reg26);
              reg35 = reg32[(2'h2):(1'h0)];
              reg36 = ((reg31[(1'h0):(1'h0)] << $unsigned(reg26)) ?
                  $unsigned(wire17[(5'h10):(2'h3)]) : ($unsigned({(~^reg30)}) ?
                      $signed($unsigned($unsigned(wire18))) : $unsigned((&$unsigned(reg35)))));
              reg37 <= (reg31 ? reg26 : $unsigned(reg31));
            end
          for (forvar38 = (1'h0); (forvar38 < (1'h1)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= (~&(reg23 << (|(7'h43))));
              reg40 <= ((+(reg34[(5'h10):(4'hb)] ?
                      reg24[(5'h10):(3'h5)] : $signed(wire18[(1'h1):(1'h0)]))) ?
                  wire16[(2'h2):(2'h2)] : ($unsigned(forvar38) ?
                      (-wire21) : ($unsigned($signed(reg31)) ^ (~(wire22 ?
                          reg35 : forvar29)))));
              reg41 <= wire19;
              reg42 = ($signed($signed($signed(reg39))) ?
                  (~^$unsigned($unsigned($signed((8'h9e))))) : {($unsigned(wire19) & {$signed(reg33),
                          (wire21 ^ forvar38)}),
                      (wire17[(4'hb):(3'h4)] <<< $signed((-(8'ha8))))});
              reg43 = "JgG0dOxXf15ygU";
            end
          if ((reg39[(3'h7):(2'h3)] ?
              (wire21[(2'h2):(1'h1)] ?
                  ($signed((8'haa)) ?
                      {reg39,
                          $unsigned(reg39)} : wire21[(3'h4):(2'h2)]) : $unsigned(((reg33 ?
                      (8'hb0) : (8'ha8)) > $signed(wire18)))) : {$unsigned(reg33),
                  wire20[(4'h9):(2'h3)]}))
            begin
              reg44 <= (((|(reg26[(3'h4):(2'h3)] ?
                      (reg24 ? (8'ha5) : wire21) : $unsigned(reg39))) ?
                  (~{$unsigned((8'ha8)),
                      (~^(8'haa))}) : $unsigned($signed("Doih6IDmV"))) >= (((^~reg23) | ((reg39 ~^ reg23) ?
                      wire19 : $unsigned(reg33))) ?
                  reg36 : $unsigned((~|reg39))));
              reg45 <= (&wire17);
              reg46 <= (7'h43);
            end
          else
            begin
              reg44 <= reg37[(2'h3):(2'h2)];
              reg45 = reg28;
              reg46 = (8'hbe);
            end
        end
      else
        begin
          reg34 = ((7'h42) ?
              (reg33 ?
                  {((|reg44) ?
                          {reg23} : (wire17 == wire19))} : ({$unsigned(forvar25),
                      reg36[(5'h10):(1'h1)]} & reg30[(4'h8):(1'h0)])) : reg26[(3'h6):(1'h1)]);
          for (forvar35 = (1'h0); (forvar35 < (3'h4)); forvar35 = (forvar35 + (1'h1)))
            begin
              reg36 = ($unsigned($unsigned(reg41)) ?
                  $unsigned($unsigned($unsigned((wire19 | forvar38)))) : (($unsigned((!(8'hbe))) ?
                          reg45 : reg23[(1'h0):(1'h0)]) ?
                      $signed($signed((~&reg40))) : (reg43[(1'h1):(1'h0)] < $signed($unsigned(reg24)))));
              reg37 <= {$unsigned("mudRMwhf8h1k")};
              reg38 <= ($signed((7'h43)) != (((&(reg24 & wire20)) ?
                  reg36 : $signed(reg35[(5'h11):(4'he)])) != {reg36[(3'h4):(3'h4)],
                  (((8'hb4) ? reg34 : (8'hb8)) ?
                      forvar25[(5'h10):(4'hd)] : (|forvar38))}));
              reg39 = reg42[(2'h2):(2'h2)];
              reg40 = wire18;
            end
          reg41 <= ($unsigned("") ?
              wire19[(4'h8):(3'h4)] : (^((^~(8'h9d)) ?
                  ($signed((8'hb2)) ?
                      {wire18} : (wire22 ?
                          (8'had) : reg43)) : ($signed(forvar25) ?
                      $unsigned((8'ha8)) : reg44[(3'h5):(3'h5)]))));
          for (forvar42 = (1'h0); (forvar42 < (1'h1)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 <= (^~({forvar42[(1'h1):(1'h0)]} ~^ $signed((&wire19))));
              reg44 <= reg43;
              reg45 = $unsigned(($unsigned($signed((reg45 ? reg40 : (8'hb9)))) ?
                  ($signed(reg38[(1'h1):(1'h1)]) ?
                      $signed((^~reg43)) : forvar35[(4'he):(1'h0)]) : (reg24 | $unsigned(wire17))));
            end
        end
      for (forvar47 = (1'h0); (forvar47 < (3'h4)); forvar47 = (forvar47 + (1'h1)))
        begin
          for (forvar48 = (1'h0); (forvar48 < (2'h3)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 = (reg36[(5'h12):(4'hb)] ?
                  (($signed($signed(reg26)) ?
                      $unsigned(reg42) : reg32) ^ reg24) : reg31);
              reg50 <= $signed(reg26);
              reg51 <= reg37[(2'h3):(2'h2)];
            end
        end
      reg52 <= forvar47;
      for (forvar53 = (1'h0); (forvar53 < (2'h3)); forvar53 = (forvar53 + (1'h1)))
        begin
          for (forvar54 = (1'h0); (forvar54 < (1'h1)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 = forvar54;
            end
        end
    end
  assign wire56 = reg52[(4'ha):(4'h9)];
  assign wire57 = {(8'haf)};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module324
#( parameter param452 = ((!(|(((7'h44) + (8'hb4)) ? {(8'had), (8'h9d)} : ((8'ha0) >= (8'hbd))))) - {((((8'hb5) ? (8'ha3) : (7'h43)) ? ((8'h9e) ? (8'ha8) : (8'ha2)) : (~&(8'hab))) >= (((8'hb0) ? (8'ha1) : (8'had)) ? (-(8'hb3)) : (~(8'hbb)))), (+((|(8'ha3)) > ((8'hb9) ? (8'hb2) : (8'hac))))}) )
(y, clk, wire328, wire327, wire326, wire325);
  output wire [(32'h5a9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire328;
  input wire signed [(4'hb):(1'h0)] wire327;
  input wire [(4'hc):(1'h0)] wire326;
  input wire [(3'h5):(1'h0)] wire325;
  reg signed [(3'h7):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar450 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg449 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg448 = (1'h0);
  reg [(5'h14):(1'h0)] forvar447 = (1'h0);
  reg [(2'h2):(1'h0)] reg446 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg445 = (1'h0);
  reg [(5'h14):(1'h0)] forvar444 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar443 = (1'h0);
  reg [(4'hb):(1'h0)] reg442 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar441 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(3'h7):(1'h0)] reg439 = (1'h0);
  reg [(5'h10):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg437 = (1'h0);
  reg [(5'h11):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg435 = (1'h0);
  reg [(4'h8):(1'h0)] reg434 = (1'h0);
  reg [(3'h6):(1'h0)] reg433 = (1'h0);
  reg [(4'hd):(1'h0)] forvar432 = (1'h0);
  reg [(5'h15):(1'h0)] reg431 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg430 = (1'h0);
  reg [(5'h15):(1'h0)] reg429 = (1'h0);
  reg [(4'hb):(1'h0)] reg428 = (1'h0);
  reg [(2'h2):(1'h0)] forvar427 = (1'h0);
  reg [(4'ha):(1'h0)] reg426 = (1'h0);
  reg [(5'h11):(1'h0)] forvar425 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg424 = (1'h0);
  reg [(5'h14):(1'h0)] reg423 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar422 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire421;
  reg signed [(3'h4):(1'h0)] reg420 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar419 = (1'h0);
  reg [(5'h15):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg414 = (1'h0);
  reg [(3'h5):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar411 = (1'h0);
  reg [(3'h5):(1'h0)] reg410 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg408 = (1'h0);
  reg [(4'hf):(1'h0)] forvar407 = (1'h0);
  reg [(4'hd):(1'h0)] reg406 = (1'h0);
  reg [(4'hf):(1'h0)] forvar405 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire404;
  wire signed [(2'h2):(1'h0)] wire403;
  reg signed [(3'h6):(1'h0)] reg402 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire401;
  reg signed [(5'h11):(1'h0)] reg400 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg399 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar397 = (1'h0);
  reg [(4'hf):(1'h0)] reg396 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg395 = (1'h0);
  reg [(5'h11):(1'h0)] forvar394 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg392 = (1'h0);
  reg [(4'ha):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg390 = (1'h0);
  reg [(5'h13):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar388 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg387 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg385 = (1'h0);
  reg [(4'hb):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar382 = (1'h0);
  reg [(4'he):(1'h0)] reg381 = (1'h0);
  reg [(5'h14):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg379 = (1'h0);
  reg [(4'hb):(1'h0)] reg378 = (1'h0);
  reg [(4'ha):(1'h0)] forvar377 = (1'h0);
  reg [(2'h2):(1'h0)] reg376 = (1'h0);
  reg [(3'h6):(1'h0)] forvar375 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar374 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg373 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire372;
  reg [(5'h15):(1'h0)] reg371 = (1'h0);
  reg [(4'hb):(1'h0)] reg370 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg368 = (1'h0);
  reg [(4'hb):(1'h0)] reg367 = (1'h0);
  reg [(2'h3):(1'h0)] reg366 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg364 = (1'h0);
  reg [(5'h12):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar362 = (1'h0);
  reg [(4'h8):(1'h0)] forvar361 = (1'h0);
  reg [(4'hf):(1'h0)] reg360 = (1'h0);
  reg [(4'hb):(1'h0)] reg359 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar358 = (1'h0);
  wire [(4'h9):(1'h0)] wire357;
  wire [(4'h8):(1'h0)] wire356;
  wire [(5'h15):(1'h0)] wire355;
  reg signed [(3'h7):(1'h0)] reg354 = (1'h0);
  reg [(3'h6):(1'h0)] reg353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg349 = (1'h0);
  reg [(4'h8):(1'h0)] reg348 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg347 = (1'h0);
  reg [(4'he):(1'h0)] reg346 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg345 = (1'h0);
  reg [(5'h14):(1'h0)] reg344 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg343 = (1'h0);
  reg signed [(4'he):(1'h0)] reg342 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg341 = (1'h0);
  reg [(3'h4):(1'h0)] reg340 = (1'h0);
  reg [(3'h4):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar335 = (1'h0);
  reg signed [(4'he):(1'h0)] reg334 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg331 = (1'h0);
  reg [(3'h6):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg337 = (1'h0);
  reg [(3'h6):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg335 = (1'h0);
  reg [(5'h15):(1'h0)] forvar334 = (1'h0);
  reg [(5'h13):(1'h0)] reg333 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg332 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar331 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg329 = (1'h0);
  assign y = {reg451,
                 forvar450,
                 reg449,
                 reg448,
                 forvar447,
                 reg446,
                 reg445,
                 forvar444,
                 forvar443,
                 reg442,
                 forvar441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 reg426,
                 forvar425,
                 reg424,
                 reg423,
                 forvar422,
                 wire421,
                 reg420,
                 forvar419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 forvar411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 forvar405,
                 wire404,
                 wire403,
                 reg402,
                 wire401,
                 reg400,
                 reg399,
                 reg398,
                 forvar397,
                 reg396,
                 reg395,
                 forvar394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 forvar388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 forvar375,
                 forvar374,
                 reg373,
                 wire372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 forvar361,
                 reg360,
                 reg359,
                 forvar358,
                 wire357,
                 wire356,
                 wire355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 forvar335,
                 reg334,
                 reg331,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 forvar334,
                 reg333,
                 reg332,
                 forvar331,
                 reg330,
                 reg329,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg329 <= (8'had);
    end
  always
    @(posedge clk) begin
      if (({((~^$signed(wire325)) ?
              wire327[(4'h9):(3'h4)] : $unsigned((wire327 > (8'hb0)))),
          (wire326 < $signed((~^wire328)))} < $signed($unsigned($signed("ncFtkNWEVL")))))
        begin
          reg330 <= (+(((~^wire328[(3'h4):(1'h1)]) && ((wire327 >= wire325) >> $signed(reg329))) ?
              reg329 : reg329[(1'h0):(1'h0)]));
          for (forvar331 = (1'h0); (forvar331 < (2'h2)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 <= (wire326 ?
                  ((~&((wire326 && wire326) ?
                          ((8'hab) ? forvar331 : wire327) : $signed(wire326))) ?
                      (($signed(wire327) ? $signed(wire328) : (&(8'ha8))) ?
                          wire327[(2'h3):(1'h1)] : "0SaC7v") : reg329[(2'h2):(1'h0)]) : (wire328[(3'h6):(1'h1)] ?
                      $signed(wire328) : (reg330[(3'h4):(2'h2)] ?
                          forvar331 : wire327[(3'h6):(3'h5)])));
              reg333 = (~$signed($signed((~^(forvar331 - reg329)))));
            end
          for (forvar334 = (1'h0); (forvar334 < (1'h0)); forvar334 = (forvar334 + (1'h1)))
            begin
              reg335 <= {forvar331};
              reg336 <= reg333;
            end
          if ($signed((+{(~|$signed(reg335))})))
            begin
              reg337 = (^$signed(wire326[(4'h8):(2'h2)]));
              reg338 <= (^(8'had));
            end
          else
            begin
              reg337 <= reg335[(5'h10):(2'h2)];
            end
        end
      else
        begin
          if ((^~{{{(wire327 ~^ reg338)}}}))
            begin
              reg330 = (8'haf);
              reg331 = $unsigned($unsigned((forvar334[(5'h12):(4'hc)] ?
                  reg335 : (!reg329[(2'h3):(1'h1)]))));
              reg332 <= $unsigned((reg333 ? "LUFbZ" : wire327));
              reg333 <= wire328;
              reg334 <= (8'hb0);
            end
          else
            begin
              reg330 = $signed($signed(((8'hb7) * reg337[(5'h14):(4'ha)])));
            end
          for (forvar335 = (1'h0); (forvar335 < (3'h4)); forvar335 = (forvar335 + (1'h1)))
            begin
              reg336 = (reg333[(3'h7):(2'h3)] && (8'haf));
              reg337 = $unsigned(($unsigned({$signed(reg335),
                  $signed(reg337)}) + {$signed(wire328)}));
              reg338 <= {reg336[(2'h2):(1'h1)]};
            end
          reg339 = $unsigned(((~((reg338 ~^ reg329) ?
              forvar334[(5'h12):(5'h10)] : "d0hNmcsx5PPCJi")) + (forvar334 ?
              $unsigned({reg337}) : (~&$signed(reg334)))));
          reg340 <= reg339[(2'h3):(1'h1)];
          if ("yVLsd181k2bI")
            begin
              reg341 = $unsigned(reg334);
            end
          else
            begin
              reg341 <= $unsigned(({"o3Mc4Kz"} || ($unsigned($signed(wire328)) - {{reg337}})));
              reg342 <= "5qyDx";
              reg343 <= ((~^reg332) ?
                  ($unsigned(((|reg341) ?
                      reg331 : $signed(reg337))) > ({(reg338 ?
                          (8'ha6) : (8'hbe)),
                      (+reg338)} && $unsigned($unsigned(reg339)))) : ((8'ha6) ?
                      (~wire327) : $unsigned(forvar331[(3'h6):(2'h3)])));
              reg344 <= ($unsigned($signed((reg337[(4'hc):(3'h7)] >= (wire327 <<< reg343)))) ?
                  (|($signed($signed(reg335)) * $signed(reg337[(5'h11):(1'h1)]))) : $unsigned(forvar331[(4'ha):(3'h5)]));
              reg345 <= (+("cVIXn5GUHDhO2w" ?
                  $signed((~&reg332)) : forvar335[(4'h9):(3'h5)]));
            end
        end
      reg346 <= $unsigned(($unsigned($unsigned(reg344[(1'h1):(1'h0)])) ?
          reg331[(4'h9):(2'h2)] : (((!reg333) ?
              (forvar335 * reg339) : $signed(reg331)) || $signed(forvar331[(2'h3):(1'h0)]))));
      if (reg336)
        begin
          reg347 = ((reg337[(5'h12):(1'h0)] == (reg332[(3'h7):(2'h2)] == (^~$unsigned(reg335)))) ?
              $signed($signed((+wire327))) : reg332[(2'h3):(1'h0)]);
          reg348 <= ((7'h41) ? wire327 : reg337);
        end
      else
        begin
          reg347 <= $unsigned(reg338[(2'h2):(1'h0)]);
          reg348 <= {(reg341 | reg335[(4'ha):(4'h8)]), reg343[(1'h0):(1'h0)]};
          if ($unsigned(reg344[(5'h14):(2'h3)]))
            begin
              reg349 = wire328;
              reg350 <= reg341[(2'h2):(1'h1)];
              reg351 <= reg338;
              reg352 <= $unsigned(reg336[(3'h6):(1'h1)]);
            end
          else
            begin
              reg349 = reg349;
              reg350 <= ((reg329[(4'hf):(2'h2)] ?
                  (-{reg329,
                      {reg349,
                          (7'h41)}}) : ((|forvar334[(5'h10):(2'h3)]) > forvar335)) && ({$signed(reg348),
                  reg341[(3'h7):(3'h5)]} ~^ $unsigned($unsigned((~reg342)))));
              reg351 = (reg351 >= (8'had));
              reg352 = (|"o9HFallJw2Zd3YoO");
            end
          reg353 <= $unsigned((^($signed($signed(forvar334)) ?
              $signed((reg352 ? reg350 : reg350)) : (reg343 ?
                  "4d" : forvar331))));
          reg354 = $signed(wire326);
        end
    end
  assign wire355 = ({(reg348 ?
                               ($signed((8'ha7)) - (reg346 ?
                                   reg333 : reg338)) : reg352)} ?
                       reg339[(2'h2):(1'h0)] : $signed($signed(((^wire328) - reg352[(2'h3):(2'h3)]))));
  assign wire356 = (((+(reg344 ? (reg334 - (8'haf)) : wire327)) ?
                           $signed(($signed(reg343) ?
                               (reg337 ?
                                   reg351 : reg337) : reg344)) : $unsigned((reg342 ?
                               $signed((7'h41)) : (forvar335 >>> forvar334)))) ?
                       $signed("") : (reg333[(3'h4):(1'h1)] ?
                           {reg335[(4'h8):(3'h7)]} : reg344[(4'hd):(3'h4)]));
  assign wire357 = forvar335;
  always
    @(posedge clk) begin
      for (forvar358 = (1'h0); (forvar358 < (1'h1)); forvar358 = (forvar358 + (1'h1)))
        begin
          if (wire325[(2'h2):(1'h1)])
            begin
              reg359 = (~&((!$unsigned((wire325 ? reg340 : reg347))) ?
                  (+(|((8'h9d) ? reg337 : forvar335))) : (wire357 ?
                      $unsigned(reg341[(4'hc):(1'h0)]) : $unsigned($unsigned(reg338)))));
            end
          else
            begin
              reg359 <= ((forvar331[(4'h8):(3'h7)] ^~ ($signed(reg342) ^ reg348[(3'h7):(3'h6)])) ?
                  $signed((~^($signed(reg345) <= reg335))) : {$signed(reg343[(1'h0):(1'h0)]),
                      {$unsigned($unsigned(reg329))}});
              reg360 = ((^~reg334[(3'h6):(2'h2)]) ?
                  $unsigned($unsigned(reg351)) : $unsigned((!$signed(reg339))));
            end
        end
      for (forvar361 = (1'h0); (forvar361 < (2'h2)); forvar361 = (forvar361 + (1'h1)))
        begin
          for (forvar362 = (1'h0); (forvar362 < (2'h2)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 = (~^$signed((-$unsigned(reg330[(4'hd):(3'h6)]))));
            end
          reg364 = ($signed((~&($signed(reg331) ?
                  {wire357, wire355} : ((8'hb5) > forvar361)))) ?
              (~^forvar331) : (|reg342[(2'h3):(2'h2)]));
          reg365 = reg350;
          if (reg342)
            begin
              reg366 = (reg345 ? reg342 : reg347);
              reg367 <= $signed({{$signed($unsigned(reg343))}});
              reg368 = (+reg333);
              reg369 = (wire325[(3'h4):(1'h0)] ?
                  reg336[(1'h1):(1'h0)] : $unsigned($unsigned({(reg332 ~^ wire355),
                      (~forvar331)})));
              reg370 <= ($unsigned($signed((|reg360[(1'h0):(1'h0)]))) >>> {reg367,
                  {($unsigned((8'hbc)) ?
                          (reg367 ? reg329 : reg346) : (reg347 <= reg339)),
                      $unsigned($signed(reg337))}});
            end
          else
            begin
              reg366 = $signed((!$unsigned(((reg344 ?
                  reg354 : reg359) >>> (reg368 ? reg347 : wire357)))));
            end
        end
      reg371 = (&$signed(forvar331[(3'h7):(3'h5)]));
    end
  assign wire372 = $signed((^~(reg366 + $signed("ThcJXM0ycZF4tRD"))));
  always
    @(posedge clk) begin
      reg373 = (~|(reg333 ?
          (^reg333[(4'hc):(3'h5)]) : (~^{$signed(reg364),
              reg344[(5'h14):(4'hc)]})));
      for (forvar374 = (1'h0); (forvar374 < (1'h0)); forvar374 = (forvar374 + (1'h1)))
        begin
          for (forvar375 = (1'h0); (forvar375 < (1'h1)); forvar375 = (forvar375 + (1'h1)))
            begin
              reg376 <= (8'ha8);
            end
          for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 <= (forvar334[(4'h9):(1'h1)] ?
                  $unsigned(reg369[(5'h14):(3'h4)]) : (~$signed(reg366[(2'h3):(1'h0)])));
              reg379 <= $unsigned($unsigned(((~|(8'ha9)) ?
                  $unsigned($unsigned(forvar358)) : wire372[(3'h4):(1'h0)])));
              reg380 <= ((!(reg350[(2'h2):(2'h2)] ?
                      "yzZcRskcH1YGa3bbB" : ((reg363 << forvar375) == reg379[(2'h3):(2'h3)]))) ?
                  (reg370[(3'h5):(2'h3)] ?
                      $unsigned((|$unsigned(wire327))) : reg338) : (((reg376 ?
                          forvar375[(1'h1):(1'h0)] : (wire326 ^ reg354)) && reg378[(1'h0):(1'h0)]) ?
                      (((wire326 > reg379) <<< ((8'haf) != forvar335)) ?
                          ((&reg338) ?
                              forvar335 : reg349) : (~|$unsigned(reg338))) : reg353));
              reg381 <= (8'had);
            end
          for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 <= ({((8'ha9) ? reg335 : (-$unsigned(reg348))), wire372} ?
                  forvar334[(5'h14):(5'h12)] : wire357);
              reg384 = (((!$signed((reg376 <= forvar374))) ^~ $unsigned(reg353)) ?
                  {$unsigned(reg331),
                      ($signed((!wire355)) ?
                          $unsigned(forvar331[(1'h0):(1'h0)]) : $unsigned((reg349 ?
                              reg366 : reg368)))} : $unsigned($unsigned({reg342[(1'h0):(1'h0)]})));
              reg385 = $signed((({reg334} != wire357) ~^ (((^reg350) <= reg343) ?
                  (reg381[(4'hc):(1'h1)] ?
                      reg338 : wire328[(3'h5):(1'h1)]) : (^$signed(reg335)))));
              reg386 = ((reg383 ?
                      (reg380 ^ $unsigned((reg341 > reg332))) : $unsigned(($signed((8'hb8)) ?
                          (reg359 ? reg341 : reg381) : reg329))) ?
                  "6vkwTZ03bu97RgmzOIik" : reg331[(3'h5):(3'h4)]);
              reg387 <= ((|$signed(reg385[(3'h6):(3'h4)])) <<< (reg359[(3'h4):(2'h3)] ?
                  (|(~&(reg381 ?
                      wire328 : reg351))) : (~|(!$unsigned(reg360)))));
            end
          for (forvar388 = (1'h0); (forvar388 < (3'h4)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 <= ($signed({$signed(reg379[(3'h7):(1'h1)]),
                  reg345}) != ((($signed(reg354) >> (reg384 ?
                      reg368 : reg349)) & $signed((~|(8'hba)))) ?
                  reg337[(5'h12):(2'h3)] : $signed((~&(wire356 ?
                      reg333 : (8'ha6))))));
              reg390 <= "Cy0ByWgsw56P5Q";
              reg391 = $signed(((|$unsigned((reg387 ? reg339 : reg390))) ?
                  $unsigned((&(-wire357))) : ($unsigned(reg364) + forvar334[(1'h1):(1'h0)])));
              reg392 = ($signed(reg384) < ((~|{(|reg338),
                  (&reg344)}) == (~(8'h9e))));
              reg393 <= $unsigned($signed((&$unsigned((^~forvar377)))));
            end
        end
      for (forvar394 = (1'h0); (forvar394 < (1'h0)); forvar394 = (forvar394 + (1'h1)))
        begin
          reg395 = reg346;
          reg396 <= wire356[(3'h5):(3'h5)];
          for (forvar397 = (1'h0); (forvar397 < (3'h4)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 = $unsigned((($signed((reg367 ?
                      reg337 : wire355)) | $signed({reg380})) ?
                  "gL5b" : $unsigned((+$unsigned((8'had))))));
            end
          reg399 = forvar394;
          reg400 <= (+$signed($signed($unsigned(forvar358))));
        end
    end
  assign wire401 = $unsigned((-reg330));
  always
    @(posedge clk) begin
      reg402 <= $unsigned((reg370 ^ (((forvar394 ^ reg360) == $signed(reg350)) ?
          $unsigned($signed(reg344)) : ($signed(reg342) ?
              $unsigned(wire372) : {forvar361}))));
    end
  assign wire403 = $unsigned({(8'had), (8'ha2)});
  assign wire404 = ((reg380 * "eehu9EBoRd9CbJ250") ?
                       ($signed((~(reg363 >> reg330))) ?
                           ((!(!reg386)) + $signed((reg399 != reg345))) : ($unsigned(reg367[(4'hb):(1'h0)]) | $unsigned(reg402))) : ({reg396} * {{{(8'ha4),
                                   reg378}},
                           {(^reg363)}}));
  always
    @(posedge clk) begin
      for (forvar405 = (1'h0); (forvar405 < (1'h0)); forvar405 = (forvar405 + (1'h1)))
        begin
          reg406 <= reg329;
          for (forvar407 = (1'h0); (forvar407 < (2'h2)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 <= reg348[(1'h1):(1'h0)];
              reg409 <= (|$unsigned((8'haf)));
              reg410 = reg333[(5'h12):(4'h9)];
            end
          for (forvar411 = (1'h0); (forvar411 < (1'h1)); forvar411 = (forvar411 + (1'h1)))
            begin
              reg412 <= reg348;
              reg413 <= (+reg336);
              reg414 = (wire403[(1'h1):(1'h1)] ?
                  $unsigned($signed($unsigned(reg337[(1'h1):(1'h1)]))) : forvar405);
              reg415 <= reg335;
            end
        end
      reg416 = $unsigned(forvar388);
      reg417 = $signed($signed($unsigned($signed((reg398 ?
          (8'h9f) : forvar394)))));
      reg418 <= reg343[(2'h2):(1'h0)];
      for (forvar419 = (1'h0); (forvar419 < (2'h2)); forvar419 = (forvar419 + (1'h1)))
        begin
          reg420 = ((~|wire404[(3'h5):(1'h0)]) ?
              ($unsigned(((reg413 ?
                      wire403 : reg385) < forvar335[(4'hd):(4'ha)])) ?
                  $signed($unsigned($signed(forvar362))) : (|reg341)) : "Z8LA7ftEs");
        end
    end
  assign wire421 = $signed((reg360 < $unsigned($unsigned($signed(wire357)))));
  always
    @(posedge clk) begin
      for (forvar422 = (1'h0); (forvar422 < (2'h2)); forvar422 = (forvar422 + (1'h1)))
        begin
          reg423 = $signed({reg406,
              $unsigned($unsigned(reg413[(2'h2):(1'h0)]))});
        end
      reg424 = reg353;
      for (forvar425 = (1'h0); (forvar425 < (2'h2)); forvar425 = (forvar425 + (1'h1)))
        begin
          reg426 <= $unsigned(reg379);
          for (forvar427 = (1'h0); (forvar427 < (3'h4)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= {$unsigned(wire355[(4'h9):(3'h7)])};
              reg429 = (($unsigned((~$signed(reg336))) ^~ (~$signed(reg386[(1'h1):(1'h0)]))) > $signed("zQTPGc6HZqvn"));
              reg430 = reg429;
              reg431 <= {($unsigned(($signed(reg416) ?
                      $unsigned(reg367) : $signed((8'hbb)))) <= $signed($unsigned($unsigned(reg369)))),
                  (forvar427[(1'h1):(1'h1)] ?
                      $signed(($signed(reg384) ?
                          "on8lm5P9GFJ4n048w" : (reg393 ?
                              (7'h40) : reg417))) : (8'hb2))};
            end
          for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= forvar361;
              reg434 <= (+{$signed($unsigned($signed(reg430)))});
              reg435 = wire327;
            end
          if (reg433[(1'h0):(1'h0)])
            begin
              reg436 = (~&($unsigned(reg379) ?
                  (forvar361[(4'h8):(1'h1)] ?
                      wire325[(3'h5):(1'h0)] : $signed($unsigned(forvar407))) : (reg351[(1'h1):(1'h0)] || (&(reg418 ?
                      reg365 : reg414)))));
              reg437 <= $signed(reg429);
              reg438 = reg399;
            end
          else
            begin
              reg436 = reg348[(4'h8):(3'h4)];
              reg437 <= wire327[(3'h7):(2'h3)];
              reg438 = forvar432[(1'h1):(1'h1)];
              reg439 <= ($unsigned(reg396[(1'h0):(1'h0)]) ?
                  reg371 : (|$unsigned(reg368)));
              reg440 <= $signed(reg341[(3'h4):(2'h2)]);
            end
          for (forvar441 = (1'h0); (forvar441 < (2'h2)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 = forvar394;
            end
        end
      for (forvar443 = (1'h0); (forvar443 < (3'h4)); forvar443 = (forvar443 + (1'h1)))
        begin
          for (forvar444 = (1'h0); (forvar444 < (2'h2)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 <= {$unsigned(reg369[(3'h4):(1'h1)])};
            end
          reg446 = $signed((7'h40));
          for (forvar447 = (1'h0); (forvar447 < (1'h0)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 <= reg370;
            end
        end
    end
  always
    @(posedge clk) begin
      reg449 = $unsigned(reg430[(3'h7):(2'h2)]);
      for (forvar450 = (1'h0); (forvar450 < (1'h1)); forvar450 = (forvar450 + (1'h1)))
        begin
          reg451 <= ($unsigned((^~forvar361[(4'h8):(3'h5)])) && (~|reg354));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module71
#( parameter param236 = (!(((8'ha6) | (((8'ha6) < (8'hb4)) ? ((7'h40) ? (8'hab) : (8'h9f)) : ((8'ha6) ? (7'h43) : (8'h9c)))) | ((((8'hbb) >>> (8'ha0)) ? ((7'h41) && (8'hbe)) : ((8'hac) >= (8'hb4))) ? (-(~(8'ha2))) : {{(7'h42), (8'hab)}, ((8'hb6) > (8'ha3))})))
, parameter param237 = (8'haa) )
(y, clk, wire76, wire75, wire74, wire73, wire72);
  output wire [(32'h763):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire76;
  input wire signed [(4'ha):(1'h0)] wire75;
  input wire signed [(5'h15):(1'h0)] wire74;
  input wire signed [(3'h5):(1'h0)] wire73;
  input wire signed [(2'h2):(1'h0)] wire72;
  wire [(4'hf):(1'h0)] wire235;
  reg [(4'hd):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg233 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar232 = (1'h0);
  reg [(4'ha):(1'h0)] reg231 = (1'h0);
  reg [(3'h7):(1'h0)] reg230 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg228 = (1'h0);
  reg [(5'h12):(1'h0)] forvar227 = (1'h0);
  reg [(2'h2):(1'h0)] reg226 = (1'h0);
  reg [(4'he):(1'h0)] reg225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg224 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg223 = (1'h0);
  reg [(3'h5):(1'h0)] reg222 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar220 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg221 = (1'h0);
  reg [(4'hd):(1'h0)] reg220 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg218 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg217 = (1'h0);
  reg signed [(4'he):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg215 = (1'h0);
  reg [(4'h9):(1'h0)] reg214 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg211 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar210 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg209 = (1'h0);
  reg [(3'h6):(1'h0)] reg208 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg207 = (1'h0);
  reg [(4'hb):(1'h0)] reg206 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar205 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg204 = (1'h0);
  reg [(3'h7):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg202 = (1'h0);
  reg [(2'h3):(1'h0)] forvar201 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar195 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(4'hc):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg197 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg196 = (1'h0);
  reg [(2'h3):(1'h0)] reg195 = (1'h0);
  reg [(3'h6):(1'h0)] reg194 = (1'h0);
  reg [(4'hd):(1'h0)] reg193 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar191 = (1'h0);
  reg [(5'h13):(1'h0)] reg190 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar188 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg186 = (1'h0);
  reg [(2'h2):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg183 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar182 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg181 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg180 = (1'h0);
  reg [(4'ha):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar178 = (1'h0);
  wire [(4'ha):(1'h0)] wire177;
  reg signed [(4'ha):(1'h0)] reg176 = (1'h0);
  reg [(4'h8):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar173 = (1'h0);
  reg [(4'hb):(1'h0)] reg172 = (1'h0);
  reg [(3'h4):(1'h0)] reg171 = (1'h0);
  reg [(4'h9):(1'h0)] reg170 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(4'he):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg166 = (1'h0);
  reg [(4'hf):(1'h0)] reg165 = (1'h0);
  reg [(3'h6):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg163 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg159 = (1'h0);
  reg [(3'h4):(1'h0)] reg158 = (1'h0);
  reg [(4'hb):(1'h0)] forvar157 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg156 = (1'h0);
  reg [(4'hd):(1'h0)] forvar155 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(4'h8):(1'h0)] forvar148 = (1'h0);
  reg [(5'h14):(1'h0)] reg154 = (1'h0);
  reg [(4'ha):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar150 = (1'h0);
  reg [(5'h12):(1'h0)] reg149 = (1'h0);
  reg [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg146 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar145 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg144 = (1'h0);
  reg [(5'h14):(1'h0)] forvar143 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire142;
  wire signed [(5'h13):(1'h0)] wire141;
  reg [(3'h6):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg139 = (1'h0);
  reg [(4'hf):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar137 = (1'h0);
  reg [(4'hd):(1'h0)] reg136 = (1'h0);
  reg [(4'ha):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg132 = (1'h0);
  reg [(2'h3):(1'h0)] reg131 = (1'h0);
  reg [(4'he):(1'h0)] forvar130 = (1'h0);
  reg [(4'h9):(1'h0)] reg129 = (1'h0);
  reg [(5'h15):(1'h0)] reg128 = (1'h0);
  reg [(4'h8):(1'h0)] forvar127 = (1'h0);
  reg [(5'h14):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar125 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire124;
  reg signed [(4'h9):(1'h0)] reg123 = (1'h0);
  reg [(4'ha):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg120 = (1'h0);
  reg [(5'h10):(1'h0)] reg119 = (1'h0);
  reg [(3'h5):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg116 = (1'h0);
  reg [(5'h12):(1'h0)] reg115 = (1'h0);
  reg [(5'h10):(1'h0)] forvar114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg111 = (1'h0);
  reg [(3'h5):(1'h0)] forvar110 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar109 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg106 = (1'h0);
  reg [(3'h7):(1'h0)] reg105 = (1'h0);
  reg [(5'h13):(1'h0)] forvar104 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar103 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire102;
  wire [(4'hd):(1'h0)] wire101;
  wire signed [(4'h9):(1'h0)] wire100;
  wire [(5'h11):(1'h0)] wire99;
  reg signed [(4'hc):(1'h0)] reg98 = (1'h0);
  reg [(4'hb):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg96 = (1'h0);
  reg [(5'h15):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar93 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg92 = (1'h0);
  reg [(3'h5):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg90 = (1'h0);
  reg [(5'h10):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg88 = (1'h0);
  reg [(5'h13):(1'h0)] forvar87 = (1'h0);
  reg [(3'h6):(1'h0)] reg86 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar85 = (1'h0);
  reg [(5'h12):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg83 = (1'h0);
  reg [(3'h7):(1'h0)] forvar82 = (1'h0);
  reg [(5'h13):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg80 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg79 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar78 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg77 = (1'h0);
  assign y = {wire235,
                 reg234,
                 reg233,
                 forvar232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 forvar227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 forvar220,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 forvar205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 forvar195,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 forvar188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 forvar182,
                 reg181,
                 reg180,
                 reg179,
                 forvar178,
                 wire177,
                 reg176,
                 reg175,
                 reg174,
                 forvar173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 forvar157,
                 reg156,
                 forvar155,
                 reg150,
                 forvar148,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 forvar150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 forvar145,
                 reg143,
                 reg144,
                 forvar143,
                 wire142,
                 wire141,
                 reg140,
                 reg139,
                 reg138,
                 forvar137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 forvar130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 forvar125,
                 wire124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 forvar114,
                 reg113,
                 reg112,
                 reg111,
                 forvar110,
                 forvar109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 forvar104,
                 forvar103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 forvar93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 forvar87,
                 reg86,
                 forvar85,
                 reg84,
                 reg83,
                 forvar82,
                 reg78,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 forvar78,
                 reg77,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg77 = wire72[(1'h0):(1'h0)];
      if ($signed(reg77))
        begin
          for (forvar78 = (1'h0); (forvar78 < (3'h4)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 <= $signed($unsigned($unsigned(($signed(reg77) <= (reg77 ?
                  wire76 : wire75)))));
              reg80 = (~^$unsigned((^~$signed((reg79 ? reg77 : wire74)))));
              reg81 <= wire74;
              reg82 = $signed($signed(({$signed(reg77),
                  (reg80 ? wire74 : reg79)} > forvar78)));
            end
        end
      else
        begin
          if (((wire76 ?
              ({wire73} ~^ reg77) : (reg82[(3'h7):(1'h1)] ^~ wire72[(1'h1):(1'h0)])) & $unsigned(forvar78[(4'h8):(3'h7)])))
            begin
              reg78 <= $unsigned($unsigned(wire75[(3'h5):(2'h2)]));
              reg79 = ((^~($unsigned(wire76) & wire73[(2'h3):(1'h1)])) - (reg78 > $signed(("uDiOYlZ1" | {reg78,
                  (8'hb8)}))));
              reg80 <= (reg82[(1'h0):(1'h0)] == {((~^reg80) ?
                      $unsigned((reg80 ? wire72 : wire72)) : (8'hb7)),
                  $unsigned(wire73[(1'h0):(1'h0)])});
              reg81 <= forvar78[(4'hc):(4'hc)];
            end
          else
            begin
              reg78 = {{"2TWY0ESo2FRAew3LP2E2"}};
            end
          for (forvar82 = (1'h0); (forvar82 < (2'h3)); forvar82 = (forvar82 + (1'h1)))
            begin
              reg83 = ($unsigned($signed(reg81[(2'h2):(1'h0)])) ?
                  reg79[(1'h0):(1'h0)] : {{$unsigned({wire76, reg81}),
                          reg81[(3'h5):(2'h2)]},
                      reg81[(3'h6):(1'h0)]});
              reg84 <= {((reg79 ?
                          ((forvar78 == wire76) ?
                              wire74 : (reg82 ?
                                  reg77 : reg79)) : (reg80[(1'h1):(1'h0)] ^ $signed(forvar78))) ?
                      $signed(wire72[(1'h0):(1'h0)]) : (({reg78,
                              wire72} >= (forvar78 > wire76)) ?
                          (^~(wire75 ? reg80 : reg78)) : ((wire76 ?
                              wire75 : reg82) | reg77[(3'h5):(3'h5)])))};
            end
          for (forvar85 = (1'h0); (forvar85 < (2'h2)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 = (-$signed($signed((^~wire72))));
            end
        end
      for (forvar87 = (1'h0); (forvar87 < (2'h3)); forvar87 = (forvar87 + (1'h1)))
        begin
          if (reg79[(2'h2):(1'h1)])
            begin
              reg88 = $signed(forvar85[(1'h1):(1'h0)]);
              reg89 <= reg77;
            end
          else
            begin
              reg88 <= (~|((((reg89 ?
                      (7'h43) : forvar78) ^ (wire74 ~^ reg79)) != (|(reg83 || reg78))) ?
                  ($unsigned($unsigned((8'ha2))) >> (((8'hb3) - (8'h9d)) || (~reg84))) : reg86));
              reg89 = ((7'h44) ?
                  $unsigned($signed(reg89[(2'h3):(1'h1)])) : wire73);
              reg90 <= ((reg89 << (+{$unsigned(wire72), (^wire72)})) ?
                  $unsigned((8'hb4)) : reg86);
              reg91 <= {reg78, wire75[(3'h4):(1'h1)]};
              reg92 <= (8'hb8);
            end
          for (forvar93 = (1'h0); (forvar93 < (1'h0)); forvar93 = (forvar93 + (1'h1)))
            begin
              reg94 = $signed($unsigned(wire76));
              reg95 = $signed($unsigned(reg82[(4'h8):(3'h7)]));
              reg96 = $unsigned($signed(({{wire75, (8'hb5)}} >= reg90)));
              reg97 <= (((forvar78 < $signed((-(8'hab)))) ?
                      reg91 : (reg83 ?
                          $unsigned((wire73 >= reg92)) : {$signed(reg96)})) ?
                  {(7'h42),
                      ($signed($signed((8'hbe))) * ({reg94,
                          (8'hbc)} >> reg86))} : reg82);
            end
        end
      reg98 = $signed($signed(($signed((~^reg84)) ?
          (reg77 ? {reg88, wire75} : reg89) : $signed((wire75 ?
              forvar85 : reg95)))));
    end
  assign wire99 = $unsigned((~^((8'hbf) ?
                      ((~&forvar78) ? reg89 : (reg89 <<< reg82)) : forvar78)));
  assign wire100 = "1EQGQTsxgrt8WlwYsOyB";
  assign wire101 = ((reg86[(1'h1):(1'h0)] ?
                           $signed(($unsigned(reg96) ?
                               (forvar82 | reg86) : $unsigned(reg89))) : $unsigned(reg88)) ?
                       ("ei9Zxs64qc7h7NkPT3K" - (&($signed(reg78) <= $signed(reg88)))) : "o");
  assign wire102 = reg91;
  always
    @(posedge clk) begin
      for (forvar103 = (1'h0); (forvar103 < (3'h4)); forvar103 = (forvar103 + (1'h1)))
        begin
          for (forvar104 = (1'h0); (forvar104 < (1'h1)); forvar104 = (forvar104 + (1'h1)))
            begin
              reg105 <= $unsigned($unsigned($signed($unsigned(((8'hbb) ^ wire72)))));
              reg106 = (reg105[(3'h5):(2'h3)] < $unsigned(reg86));
            end
          reg107 = (8'hb5);
        end
      reg108 <= (((wire99 | reg78) << ($signed(reg79[(1'h0):(1'h0)]) >>> ($unsigned(reg79) ?
              $signed(reg96) : reg80))) ?
          reg90[(1'h1):(1'h0)] : ((((^~wire102) < (forvar87 & (8'ha3))) ?
              $unsigned(reg89[(3'h5):(2'h2)]) : reg88) ^~ {forvar78[(1'h0):(1'h0)],
              wire74}));
      for (forvar109 = (1'h0); (forvar109 < (1'h0)); forvar109 = (forvar109 + (1'h1)))
        begin
          for (forvar110 = (1'h0); (forvar110 < (2'h2)); forvar110 = (forvar110 + (1'h1)))
            begin
              reg111 <= {wire76};
              reg112 <= (reg82[(3'h4):(1'h1)] >> reg92[(4'hc):(3'h7)]);
            end
          reg113 = $unsigned({reg94, reg111});
          for (forvar114 = (1'h0); (forvar114 < (3'h4)); forvar114 = (forvar114 + (1'h1)))
            begin
              reg115 <= (|$unsigned((~|((forvar103 ?
                  wire99 : wire75) | ((8'hb0) ? reg88 : reg81)))));
              reg116 <= reg98;
              reg117 <= "o0";
              reg118 = $unsigned(((+reg86) ?
                  ((~{reg80, wire100}) ?
                      reg97 : $unsigned(((8'ha4) ?
                          wire74 : reg112))) : $unsigned($unsigned("cda"))));
            end
          if ({$signed(reg106),
              (($unsigned((forvar109 ^~ forvar103)) ?
                      $unsigned(reg80[(1'h0):(1'h0)]) : $unsigned($unsigned(reg115))) ?
                  (~&(~&(reg79 ? forvar104 : reg107))) : reg84)})
            begin
              reg119 = (~&wire100);
              reg120 = (($unsigned(forvar104[(3'h5):(1'h1)]) >= $signed($unsigned(forvar110))) >= $signed(reg116[(3'h6):(3'h5)]));
              reg121 = {$signed((8'hab)), $unsigned(reg95)};
              reg122 <= $unsigned(((($unsigned((8'hb2)) ?
                  (forvar103 ?
                      reg107 : (7'h40)) : {reg113}) < reg94) | (8'haf)));
              reg123 = (reg92[(4'h8):(1'h1)] << (~^(forvar78 ?
                  forvar103 : $signed(((8'ha4) >> reg89)))));
            end
          else
            begin
              reg119 = $signed((^~$signed(forvar87[(2'h2):(1'h0)])));
              reg120 = forvar110[(3'h5):(3'h5)];
            end
        end
    end
  assign wire124 = $signed($signed((!$signed((!(8'ha4))))));
  always
    @(posedge clk) begin
      for (forvar125 = (1'h0); (forvar125 < (2'h3)); forvar125 = (forvar125 + (1'h1)))
        begin
          reg126 <= wire124;
          for (forvar127 = (1'h0); (forvar127 < (2'h2)); forvar127 = (forvar127 + (1'h1)))
            begin
              reg128 <= $signed($unsigned($unsigned($unsigned(reg117[(5'h12):(2'h2)]))));
              reg129 <= reg115[(4'hf):(4'h9)];
            end
        end
      for (forvar130 = (1'h0); (forvar130 < (1'h0)); forvar130 = (forvar130 + (1'h1)))
        begin
          if ($unsigned(reg119))
            begin
              reg131 <= reg112[(4'hd):(3'h7)];
              reg132 <= (!(reg91[(1'h0):(1'h0)] & $signed(forvar78)));
              reg133 <= reg91[(2'h3):(1'h1)];
            end
          else
            begin
              reg131 = (~^reg122[(4'ha):(4'h8)]);
              reg132 <= ($signed((8'ha3)) ?
                  reg91 : (reg89[(1'h1):(1'h0)] && {($signed(reg117) << (~wire72)),
                      reg128}));
              reg133 <= $signed({(+((|forvar78) ~^ (reg84 ? reg91 : wire124))),
                  $signed(reg123)});
              reg134 <= reg111[(3'h5):(1'h0)];
              reg135 <= ($unsigned(reg116) | forvar78);
            end
          reg136 = ((^(+($signed((7'h41)) ? {reg132, reg115} : reg123))) ?
              ($signed(({(7'h44), reg82} ?
                  (forvar127 - reg108) : (reg133 ?
                      reg135 : forvar130))) ^ (reg90[(1'h0):(1'h0)] ?
                  forvar104[(3'h5):(3'h5)] : reg98)) : reg94[(2'h3):(1'h1)]);
        end
      for (forvar137 = (1'h0); (forvar137 < (2'h3)); forvar137 = (forvar137 + (1'h1)))
        begin
          reg138 <= wire74[(1'h1):(1'h1)];
          reg139 = $signed((~|$signed(reg120)));
        end
      reg140 <= {{($signed({forvar130, (8'hbd)}) ?
                  (-(wire74 ? reg134 : forvar82)) : $signed($signed(reg139))),
              ({(-forvar93), (reg86 ? (8'h9e) : reg106)} ?
                  reg121[(1'h1):(1'h1)] : reg94[(1'h1):(1'h1)])}};
    end
  assign wire141 = $signed((forvar110 != reg88));
  assign wire142 = (($unsigned((&reg138[(4'he):(3'h5)])) ?
                           (((~&reg113) ?
                               (|forvar127) : $signed(reg119)) == $unsigned($unsigned(reg122))) : (^~reg92)) ?
                       reg95[(5'h10):(1'h0)] : forvar93[(4'hd):(4'h8)]);
  always
    @(posedge clk) begin
      if (forvar127[(2'h3):(1'h1)])
        begin
          for (forvar143 = (1'h0); (forvar143 < (2'h2)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 <= $unsigned(($unsigned($unsigned((reg80 <<< reg140))) || $signed($unsigned((!reg106)))));
            end
        end
      else
        begin
          reg143 <= "r6i";
          reg144 <= ($unsigned($unsigned(reg78)) ?
              $signed({(^~{reg95, forvar130})}) : (($unsigned((reg78 ?
                      forvar109 : reg128)) > $signed((wire124 <= reg80))) ?
                  ((7'h43) ?
                      $signed((reg98 ?
                          reg129 : reg95)) : $unsigned(reg119)) : (+((reg120 == (7'h43)) <<< ((8'h9e) > forvar130)))));
        end
      if ($unsigned((((~&$unsigned((8'hb1))) ?
          forvar127[(2'h2):(1'h1)] : (~&reg133)) ^ (reg115 == "mafT"))))
        begin
          for (forvar145 = (1'h0); (forvar145 < (3'h4)); forvar145 = (forvar145 + (1'h1)))
            begin
              reg146 <= reg98[(4'h9):(4'h9)];
              reg147 <= (((~^$unsigned((reg95 ? wire76 : wire142))) ?
                      (~$signed(reg97[(4'h8):(3'h4)])) : $signed(reg86[(3'h4):(3'h4)])) ?
                  ($signed(($unsigned(wire73) ?
                          (^reg118) : $unsigned(reg138))) ?
                      (~|forvar127) : reg96) : ((wire73 != reg115) & (-$unsigned({reg113,
                      reg95}))));
              reg148 <= reg90;
              reg149 <= $signed((((^~(8'hbf)) ?
                  $signed({forvar78}) : (reg113[(4'hc):(1'h0)] < $unsigned(forvar87))) | ($unsigned(reg106[(2'h3):(2'h3)]) && forvar110[(3'h5):(1'h0)])));
            end
          for (forvar150 = (1'h0); (forvar150 < (1'h0)); forvar150 = (forvar150 + (1'h1)))
            begin
              reg151 = reg116;
              reg152 = ((^(((!reg80) ?
                  forvar127[(1'h1):(1'h1)] : "LAwb4cunOGZoP2sYve8t") << reg113)) == $unsigned($unsigned($unsigned((reg147 > reg115)))));
              reg153 <= (8'had);
            end
          reg154 = (^~(!$unsigned(reg144)));
        end
      else
        begin
          for (forvar145 = (1'h0); (forvar145 < (1'h0)); forvar145 = (forvar145 + (1'h1)))
            begin
              reg146 = (forvar145[(1'h0):(1'h0)] <= ((7'h41) ?
                  $unsigned(wire102[(1'h1):(1'h0)]) : (reg94 ?
                      (8'hbd) : ($signed(reg88) & $signed(reg129)))));
              reg147 = reg90;
            end
          for (forvar148 = (1'h0); (forvar148 < (1'h0)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 <= "IWiBdmh";
              reg150 <= $signed(reg81);
              reg151 = (reg78[(3'h6):(1'h1)] ?
                  (reg82[(3'h4):(3'h4)] <= $unsigned(($unsigned(forvar78) <<< (wire76 >>> reg148)))) : (|($unsigned({reg96}) ?
                      $signed(forvar82[(3'h6):(3'h5)]) : reg115[(3'h4):(2'h2)])));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar155 = (1'h0); (forvar155 < (2'h2)); forvar155 = (forvar155 + (1'h1)))
        begin
          reg156 = $unsigned("U82WO");
          for (forvar157 = (1'h0); (forvar157 < (2'h2)); forvar157 = (forvar157 + (1'h1)))
            begin
              reg158 <= reg113;
              reg159 <= reg108[(2'h3):(2'h3)];
              reg160 = $unsigned({(|(reg140[(2'h2):(2'h2)] * $unsigned(forvar127)))});
              reg161 = (reg160 ?
                  $signed(((forvar109[(4'h9):(3'h7)] >>> $signed(forvar114)) ?
                      ((|forvar127) ?
                          {forvar155} : reg146) : (~$signed(reg159)))) : $signed(($signed((~(8'hb1))) ?
                      ({reg136, reg106} ?
                          (wire142 ?
                              forvar127 : forvar143) : reg97) : (reg83[(4'hb):(4'h8)] ?
                          (reg115 ^ reg84) : (reg117 | reg113)))));
              reg162 = (&reg140);
            end
          reg163 <= (|($unsigned((+(forvar150 ? reg135 : reg89))) ?
              {reg86[(1'h0):(1'h0)], $signed((|reg111))} : $unsigned((((8'ha2) ?
                      wire99 : reg158) ?
                  (+reg139) : $signed(forvar104)))));
        end
    end
  always
    @(posedge clk) begin
      reg164 <= (7'h42);
      if (reg115)
        begin
          reg165 <= $signed(reg95[(4'hf):(1'h0)]);
          reg166 = (reg161 ^ reg94);
          if ({reg90[(4'h9):(3'h6)], reg129[(4'h9):(3'h4)]})
            begin
              reg167 = reg139;
              reg168 <= $unsigned(reg163);
              reg169 <= $signed($signed((("98zbJr1kYeE4QY" ?
                  ((8'ha5) * reg97) : (+reg94)) || (forvar137[(3'h5):(1'h0)] != (reg134 ^~ (8'hbe))))));
              reg170 <= $signed($unsigned($unsigned(((-reg79) >= $unsigned(reg164)))));
              reg171 <= $signed(forvar110[(3'h5):(1'h1)]);
            end
          else
            begin
              reg167 <= wire102[(2'h2):(1'h1)];
            end
          reg172 <= (-((~$signed($unsigned(reg120))) ?
              {($unsigned(wire102) & (wire72 + reg150))} : {(+$unsigned(reg122)),
                  ({reg164, (8'hb5)} ? reg113 : (forvar103 ^ reg106))}));
          for (forvar173 = (1'h0); (forvar173 < (2'h2)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 <= ($unsigned($unsigned(reg170[(2'h3):(2'h2)])) ^~ reg151);
              reg175 <= (wire99 > $unsigned((^reg169)));
              reg176 <= (($unsigned($unsigned($signed(reg81))) >>> $unsigned(forvar82[(3'h5):(1'h0)])) ?
                  $signed((~|reg123)) : "gNUW2JWhpZSgXV");
            end
        end
      else
        begin
          if ($signed(((~$signed(forvar127)) ?
              ((&$unsigned(reg162)) ^~ (reg165[(4'h9):(1'h1)] ?
                  wire141[(4'hf):(4'h9)] : ((8'hb4) ~^ reg119))) : (!reg120))))
            begin
              reg165 = $unsigned((($signed(reg152) <= $unsigned($signed(reg91))) ?
                  forvar82[(1'h1):(1'h0)] : (&(~&$signed(reg161)))));
              reg166 = (((!$signed((!reg120))) ?
                  $unsigned((~^reg138)) : $signed((wire72[(1'h1):(1'h0)] ~^ (reg133 ?
                      wire75 : forvar114)))) >> reg107[(3'h4):(3'h4)]);
              reg167 = ($signed((+reg86)) ?
                  $unsigned((-(~^(^~forvar137)))) : ($unsigned(($unsigned(reg121) | $signed(reg146))) ?
                      reg170[(2'h3):(2'h3)] : {$unsigned(((8'ha1) ?
                              forvar78 : reg78)),
                          (-reg161)}));
            end
          else
            begin
              reg165 <= (&reg82[(1'h0):(1'h0)]);
              reg166 <= {{(~&$unsigned((forvar150 + (7'h44)))),
                      (((|reg106) ?
                          reg94[(2'h3):(2'h3)] : reg168[(2'h2):(1'h1)]) && wire74[(3'h4):(1'h1)])},
                  (+$signed((|{(8'ha1)})))};
            end
          reg168 <= reg135[(1'h0):(1'h0)];
        end
    end
  assign wire177 = (reg166 <= reg168);
  always
    @(posedge clk) begin
      for (forvar178 = (1'h0); (forvar178 < (1'h0)); forvar178 = (forvar178 + (1'h1)))
        begin
          if ({{($unsigned(((8'ha8) != wire99)) < (reg118[(2'h2):(1'h0)] ?
                      (8'hb3) : {reg122, reg171}))},
              ($signed($unsigned($signed(reg132))) || ({$unsigned(reg116),
                  $unsigned(reg118)} <= wire75))})
            begin
              reg179 <= $signed("D3MQUly");
              reg180 <= $unsigned($unsigned($signed(((+reg83) | (reg151 ?
                  reg78 : reg176)))));
              reg181 = (forvar103 ?
                  reg167[(3'h7):(1'h1)] : ((~&(+(|wire100))) | $signed(((reg147 ?
                      (8'hac) : reg135) | {reg90}))));
            end
          else
            begin
              reg179 <= wire177[(3'h5):(1'h0)];
            end
          for (forvar182 = (1'h0); (forvar182 < (2'h3)); forvar182 = (forvar182 + (1'h1)))
            begin
              reg183 = (((-((~|forvar130) || (reg106 <<< reg97))) ?
                      $unsigned(($signed((7'h43)) - ((8'hbb) ?
                          (8'ha6) : reg96))) : (reg166[(3'h5):(3'h4)] >> (~^{forvar78,
                          reg90}))) ?
                  (^~$unsigned(reg117)) : "Wf0pD81Xe1FSg");
              reg184 <= $signed($unsigned(forvar114[(4'hf):(4'hf)]));
              reg185 = forvar173;
              reg186 = reg98[(2'h3):(1'h1)];
              reg187 <= {$signed(((reg113[(3'h4):(2'h2)] ?
                          (!reg113) : {reg112, wire99}) ?
                      wire74 : forvar104)),
                  $unsigned({reg143[(3'h4):(2'h3)]})};
            end
          for (forvar188 = (1'h0); (forvar188 < (3'h4)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= $unsigned({reg135[(2'h3):(1'h1)]});
              reg190 = $signed((8'ha7));
            end
        end
      if ((((~&{(reg160 ? reg122 : reg129)}) ?
          reg105 : (reg123 + {(^~(8'hbf)),
              ((8'ha5) ?
                  (7'h43) : reg174)})) && $signed({$unsigned($unsigned(reg156))})))
        begin
          for (forvar191 = (1'h0); (forvar191 < (1'h0)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= $unsigned(((reg107 ?
                  $signed($signed(forvar182)) : ({(8'hb2),
                      reg107} > reg135)) >= ((reg184 | (forvar130 + reg144)) ?
                  (~^forvar127[(3'h6):(2'h3)]) : (forvar85 ?
                      wire76[(4'h8):(2'h3)] : $unsigned(reg147)))));
              reg193 <= $unsigned((~^reg167));
              reg194 <= wire142;
              reg195 <= ((~&(reg126 ~^ (forvar145 ?
                  (reg149 > reg153) : $unsigned(forvar145)))) != ($signed(($unsigned(reg121) ?
                  (^reg126) : (|forvar188))) >> $signed($unsigned(((7'h43) ?
                  reg146 : forvar157)))));
            end
          reg196 <= (($unsigned((reg194 ?
                  reg186[(3'h4):(3'h4)] : reg190)) + (reg180 == ($unsigned(forvar104) ?
                  (8'hbe) : (reg117 ? (8'had) : forvar130)))) ?
              reg83 : {$signed("RqdvOkEvQXcT"), reg161[(4'ha):(1'h1)]});
          reg197 <= $signed((reg78 ?
              $unsigned(reg94) : (((reg123 ? (8'ha2) : wire76) ?
                  reg161[(4'hb):(3'h6)] : reg89[(3'h6):(3'h4)]) ~^ $signed($unsigned(reg144)))));
          if (reg164[(3'h5):(1'h0)])
            begin
              reg198 <= reg175[(2'h3):(2'h3)];
              reg199 <= (&$signed(reg179[(3'h5):(2'h3)]));
              reg200 <= (reg77[(2'h3):(2'h3)] - $signed($signed(((reg116 ?
                      (8'hbd) : reg185) ?
                  reg94 : $signed(forvar148)))));
              reg201 <= $unsigned("GU3Pf3hfLQsv0dOy");
            end
          else
            begin
              reg198 <= ($signed(forvar145[(3'h7):(3'h4)]) ~^ (!$signed(reg186[(3'h5):(1'h0)])));
              reg199 <= {(~^(+$signed(reg181[(4'he):(2'h3)]))),
                  ((~|$signed((reg153 ? reg79 : reg94))) ?
                      (forvar103 >>> (!(reg126 ?
                          reg111 : reg150))) : (~^forvar182))};
              reg200 <= (8'hb2);
            end
        end
      else
        begin
          for (forvar191 = (1'h0); (forvar191 < (1'h0)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= reg79;
              reg193 = (^~$signed((8'hae)));
              reg194 = (8'hb9);
            end
          for (forvar195 = (1'h0); (forvar195 < (2'h3)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 <= (^~($signed({wire74, (~^reg154)}) ?
                  {(reg106[(2'h3):(1'h1)] ?
                          $unsigned((8'ha6)) : $signed(reg161))} : reg84));
              reg197 = reg139[(1'h1):(1'h0)];
              reg198 <= {(+"DD0PLvLVCAf1Zc")};
              reg199 <= wire102[(1'h1):(1'h1)];
              reg200 <= {(|wire141)};
            end
          for (forvar201 = (1'h0); (forvar201 < (2'h2)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 <= (($signed($signed($unsigned(forvar191))) ^~ $signed("tZXQ5N29in7Y1emzd")) ?
                  (^{$signed(reg121)}) : $unsigned(reg117[(3'h6):(3'h4)]));
              reg203 = $unsigned(({$signed(((7'h40) < reg165)),
                  (~|reg77[(3'h5):(2'h2)])} != {(-((8'haa) ?
                      reg128 : forvar103)),
                  $unsigned($unsigned(reg190))}));
              reg204 = $signed(((({(8'hae)} ?
                      (+reg136) : (reg149 ? reg175 : wire99)) ?
                  $unsigned($signed(reg91)) : $signed((reg120 ?
                      forvar109 : reg83))) | (({reg186} == $signed(reg175)) << ("uMI4D3ECDPlN9qufxWo" <= ((8'ha2) ?
                  forvar145 : reg196)))));
            end
          for (forvar205 = (1'h0); (forvar205 < (2'h3)); forvar205 = (forvar205 + (1'h1)))
            begin
              reg206 <= $unsigned("ER");
              reg207 <= (reg174[(3'h5):(2'h3)] + $signed($signed(wire74)));
              reg208 <= {(-{((reg121 - forvar93) ^ reg92[(4'ha):(4'h9)])}),
                  $unsigned(($signed((wire124 || reg126)) ?
                      reg86 : {forvar137, {reg95}}))};
              reg209 <= $unsigned($signed($unsigned({(reg129 <<< (8'ha9)),
                  (reg190 ? reg150 : reg92)})));
            end
        end
      for (forvar210 = (1'h0); (forvar210 < (1'h0)); forvar210 = (forvar210 + (1'h1)))
        begin
          if (($unsigned((^({forvar195, wire102} ?
                  ((8'ha3) ? reg184 : wire101) : (reg89 == reg187)))) ?
              reg92[(3'h5):(2'h2)] : (!($signed((reg154 && reg158)) ?
                  ($unsigned(reg129) <= (|(8'hbd))) : $unsigned(reg83[(2'h2):(1'h1)])))))
            begin
              reg211 = $signed(reg81[(1'h1):(1'h1)]);
              reg212 = ((8'ha9) || forvar191);
              reg213 = reg105;
              reg214 = "0Kztim";
            end
          else
            begin
              reg211 <= {$unsigned({$signed($signed(reg105)),
                      {{reg190, reg169}, (reg89 ? forvar191 : reg174)}})};
              reg212 <= (reg97[(2'h2):(2'h2)] >= forvar130[(3'h7):(2'h3)]);
            end
          if ($signed((~reg147[(3'h7):(2'h2)])))
            begin
              reg215 = {(+(~|$signed($signed(reg176)))),
                  (&$signed({(7'h44), (reg116 ^~ reg116)}))};
              reg216 = ($signed(wire177) ?
                  $signed((forvar125[(1'h0):(1'h0)] ?
                      $signed(forvar93[(4'h9):(3'h7)]) : ((^~(7'h44)) * {reg214,
                          reg193}))) : {(($unsigned(reg211) & (^reg135)) ?
                          {(reg186 ? forvar125 : forvar78),
                              "Od1B"} : $signed(forvar103[(2'h2):(1'h1)]))});
              reg217 <= ((~$unsigned($unsigned(reg166[(2'h2):(2'h2)]))) | (reg108[(4'h9):(3'h5)] ?
                  (($signed(forvar157) ?
                          forvar155[(4'ha):(1'h0)] : (~^wire142)) ?
                      (~reg98[(2'h2):(1'h1)]) : $signed((reg206 ?
                          reg112 : (8'hbb)))) : ((8'hb0) | ({reg96} ?
                      "" : forvar103[(1'h1):(1'h0)]))));
              reg218 = ($unsigned(reg207[(4'h8):(3'h4)]) ?
                  reg164 : $unsigned($unsigned($signed((!reg147)))));
              reg219 <= reg175;
            end
          else
            begin
              reg215 = $signed(reg95);
            end
        end
      if ((({((reg200 ? reg84 : reg148) ?
                  (reg119 ^~ reg143) : $unsigned(reg172))} <<< (forvar173 ?
              {(reg181 ? reg208 : (8'h9e)),
                  $signed(forvar210)} : reg134[(4'hb):(4'h9)])) ?
          reg139[(1'h1):(1'h1)] : (!$signed(reg165))))
        begin
          reg220 <= {(~reg128), (8'hb9)};
          reg221 <= reg161[(4'hb):(2'h2)];
        end
      else
        begin
          for (forvar220 = (1'h0); (forvar220 < (2'h2)); forvar220 = (forvar220 + (1'h1)))
            begin
              reg221 = (~|$signed((reg186 ?
                  (~^(~&reg195)) : (((8'hb1) || reg134) <<< forvar205[(4'h9):(3'h4)]))));
              reg222 = ($signed({((forvar173 << reg111) ?
                      ((8'ha8) ? reg221 : forvar109) : $signed((7'h44))),
                  reg185[(1'h0):(1'h0)]}) && reg90[(5'h10):(1'h1)]);
              reg223 = (($signed(((forvar103 << reg200) ~^ $unsigned(reg174))) ?
                  reg82 : (reg82 ? reg123 : (8'had))) | (^~{(forvar188 ?
                      (reg143 >>> reg81) : forvar87[(4'hc):(1'h1)]),
                  reg136[(2'h2):(2'h2)]}));
              reg224 <= ($signed(reg185[(2'h2):(1'h0)]) ?
                  ((($signed(reg144) || $signed((8'hbc))) >= (8'hb1)) * reg160) : ((8'h9d) <<< (8'ha6)));
            end
          reg225 <= ({({(forvar150 <= wire142), (forvar201 << reg159)} ?
                  reg119[(4'hf):(4'h9)] : $signed(((8'hbe) <<< (7'h43))))} == $unsigned(reg78[(4'h9):(4'h8)]));
          reg226 = wire76[(3'h7):(1'h1)];
          for (forvar227 = (1'h0); (forvar227 < (3'h4)); forvar227 = (forvar227 + (1'h1)))
            begin
              reg228 = reg138[(2'h3):(1'h1)];
              reg229 = {reg197};
              reg230 <= ((|(reg221[(4'hf):(2'h3)] + reg204[(2'h3):(1'h0)])) ^~ reg152[(4'h8):(3'h5)]);
              reg231 = reg217[(1'h1):(1'h0)];
            end
          for (forvar232 = (1'h0); (forvar232 < (2'h2)); forvar232 = (forvar232 + (1'h1)))
            begin
              reg233 <= (!(((^reg214) << (reg194 - reg156)) ?
                  (((reg92 ? reg151 : (8'hb3)) ?
                          (~^reg116) : (wire100 >> reg131)) ?
                      $unsigned(wire124) : wire74) : {{(reg151 ?
                              (8'hbe) : reg195)},
                      (~^{reg176})}));
            end
        end
      reg234 <= $unsigned($unsigned($unsigned({(forvar201 ? reg123 : reg107),
          (reg208 ? reg77 : (8'hbd))})));
    end
  assign wire235 = $signed("8r95M2aDNO1JHV2KfH4");
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'heb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire0;
  input wire [(4'hf):(1'h0)] wire1;
  input wire signed [(4'hb):(1'h0)] wire2;
  input wire signed [(5'h11):(1'h0)] wire3;
  wire [(2'h2):(1'h0)] wire725;
  wire signed [(5'h10):(1'h0)] wire714;
  wire [(4'h8):(1'h0)] wire713;
  wire signed [(4'he):(1'h0)] wire711;
  wire [(4'he):(1'h0)] wire710;
  reg signed [(4'hf):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar707 = (1'h0);
  reg [(5'h12):(1'h0)] reg706 = (1'h0);
  reg [(4'hd):(1'h0)] reg705 = (1'h0);
  reg [(3'h4):(1'h0)] reg704 = (1'h0);
  wire signed [(4'he):(1'h0)] wire699;
  wire signed [(5'h15):(1'h0)] wire701;
  wire [(5'h10):(1'h0)] wire702;
  wire signed [(5'h10):(1'h0)] wire716;
  wire [(3'h7):(1'h0)] wire718;
  reg [(3'h6):(1'h0)] reg720 = (1'h0);
  wire [(2'h3):(1'h0)] wire721;
  wire signed [(3'h5):(1'h0)] wire722;
  wire [(4'h8):(1'h0)] wire723;
  assign y = {wire725,
                 wire714,
                 wire713,
                 wire711,
                 wire710,
                 reg709,
                 reg708,
                 forvar707,
                 reg706,
                 reg705,
                 reg704,
                 wire699,
                 wire701,
                 wire702,
                 wire716,
                 wire718,
                 reg720,
                 wire721,
                 wire722,
                 wire723,
                 (1'h0)};
  module4 modinst700 (.y(wire699), .wire5(wire1), .wire7(wire0), .wire6(wire2), .wire9((7'h43)), .clk(clk), .wire8(wire3));
  assign wire701 = wire699;
  module4 modinst703 (wire702, clk, wire699, wire1, wire0, wire701, wire2);
  always
    @(posedge clk) begin
      reg704 <= wire1;
      reg705 <= reg704[(3'h4):(2'h3)];
      reg706 = wire1[(4'he):(2'h2)];
      for (forvar707 = (1'h0); (forvar707 < (1'h0)); forvar707 = (forvar707 + (1'h1)))
        begin
          reg708 <= wire0[(4'h8):(1'h1)];
          reg709 = (8'hb5);
        end
    end
  assign wire710 = ((8'hbe) ?
                       ($unsigned(reg704[(3'h4):(1'h1)]) >>> "KWhDo3KQ") : (8'ha2));
  module565 modinst712 (.wire566(wire710), .wire568(reg709), .wire569(wire702), .y(wire711), .clk(clk), .wire567(wire701));
  assign wire713 = $unsigned($unsigned(($signed((8'h9f)) ?
                       ($signed((8'h9d)) >> (reg705 <= wire699)) : $unsigned((forvar707 ?
                           wire3 : (8'ha7))))));
  module4 modinst715 (.wire7(forvar707), .wire6(wire701), .y(wire714), .clk(clk), .wire9(wire1), .wire8(reg705), .wire5(wire710));
  module517 modinst717 (wire716, clk, reg706, wire714, wire711, forvar707);
  module517 modinst719 (wire718, clk, wire711, reg708, wire710, wire702);
  always
    @(posedge clk) begin
      reg720 <= wire2[(2'h3):(1'h1)];
    end
  assign wire721 = (!{$unsigned(forvar707)});
  assign wire722 = wire714[(1'h1):(1'h0)];
  module270 modinst724 (.clk(clk), .wire274(wire1), .y(wire723), .wire273(wire701), .wire272(wire711), .wire275(wire699), .wire271(wire0));
  assign wire725 = $unsigned("gA7rf5N");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4  (y, clk, wire5, wire6, wire7, wire8, wire9);
  output wire [(32'h47c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire5;
  input wire signed [(2'h3):(1'h0)] wire6;
  input wire [(4'hd):(1'h0)] wire7;
  input wire signed [(4'hd):(1'h0)] wire8;
  input wire [(4'ha):(1'h0)] wire9;
  wire signed [(4'hf):(1'h0)] wire698;
  wire signed [(3'h5):(1'h0)] wire10;
  reg signed [(5'h13):(1'h0)] forvar11 = (1'h0);
  reg [(5'h14):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg14 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg15 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg17 = (1'h0);
  reg [(3'h4):(1'h0)] reg18 = (1'h0);
  reg [(4'hd):(1'h0)] forvar19 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar20 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg21 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg22 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg23 = (1'h0);
  reg [(2'h3):(1'h0)] reg24 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg25 = (1'h0);
  reg [(2'h2):(1'h0)] forvar26 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg27 = (1'h0);
  reg [(5'h10):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar27 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg29 = (1'h0);
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar32 = (1'h0);
  reg [(4'hd):(1'h0)] reg33 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg34 = (1'h0);
  reg [(2'h2):(1'h0)] reg35 = (1'h0);
  reg [(3'h6):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg37 = (1'h0);
  reg [(3'h4):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg39 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg40 = (1'h0);
  reg [(4'hd):(1'h0)] reg41 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg42 = (1'h0);
  reg [(5'h15):(1'h0)] forvar38 = (1'h0);
  reg [(4'hd):(1'h0)] forvar43 = (1'h0);
  reg [(3'h6):(1'h0)] forvar44 = (1'h0);
  reg [(3'h7):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg47 = (1'h0);
  wire [(4'h8):(1'h0)] wire48;
  reg signed [(2'h2):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg50 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire51;
  reg [(5'h12):(1'h0)] reg52 = (1'h0);
  reg [(4'hf):(1'h0)] forvar53 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg54 = (1'h0);
  reg [(5'h12):(1'h0)] reg55 = (1'h0);
  reg [(4'hc):(1'h0)] reg56 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg57 = (1'h0);
  reg [(3'h4):(1'h0)] forvar58 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg60 = (1'h0);
  reg [(5'h12):(1'h0)] reg61 = (1'h0);
  reg [(4'h8):(1'h0)] reg62 = (1'h0);
  reg [(3'h5):(1'h0)] forvar63 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg64 = (1'h0);
  reg [(5'h15):(1'h0)] reg65 = (1'h0);
  reg [(4'hc):(1'h0)] forvar66 = (1'h0);
  reg [(4'h9):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg68 = (1'h0);
  reg [(5'h10):(1'h0)] reg69 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg70 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar71 = (1'h0);
  reg [(3'h5):(1'h0)] reg72 = (1'h0);
  reg [(5'h13):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg74 = (1'h0);
  reg [(5'h11):(1'h0)] forvar75 = (1'h0);
  reg [(4'he):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg78 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire79;
  reg signed [(5'h14):(1'h0)] forvar80 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg84 = (1'h0);
  reg [(2'h3):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar86 = (1'h0);
  reg [(5'h12):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg88 = (1'h0);
  reg [(5'h12):(1'h0)] forvar89 = (1'h0);
  reg [(4'h9):(1'h0)] forvar90 = (1'h0);
  reg [(4'h8):(1'h0)] reg91 = (1'h0);
  reg [(4'he):(1'h0)] reg92 = (1'h0);
  reg [(5'h14):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg94 = (1'h0);
  reg [(4'hc):(1'h0)] reg95 = (1'h0);
  reg [(3'h5):(1'h0)] reg96 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar97 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg98 = (1'h0);
  reg [(3'h7):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg102 = (1'h0);
  reg [(4'hc):(1'h0)] reg103 = (1'h0);
  wire [(4'h9):(1'h0)] wire694;
  wire signed [(4'h8):(1'h0)] wire696;
  assign y = {wire698,
                 wire10,
                 forvar11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 forvar19,
                 forvar20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 forvar26,
                 reg27,
                 reg28,
                 reg26,
                 forvar27,
                 reg29,
                 reg30,
                 reg31,
                 forvar32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 forvar38,
                 forvar43,
                 forvar44,
                 reg45,
                 reg46,
                 reg47,
                 wire48,
                 reg49,
                 reg50,
                 wire51,
                 reg52,
                 forvar53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 forvar58,
                 reg59,
                 reg60,
                 reg61,
                 reg62,
                 forvar63,
                 reg64,
                 reg65,
                 forvar66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 forvar71,
                 reg72,
                 reg73,
                 reg74,
                 forvar75,
                 reg76,
                 reg77,
                 reg78,
                 wire79,
                 forvar80,
                 forvar81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 forvar86,
                 reg87,
                 reg88,
                 forvar89,
                 forvar90,
                 reg91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 forvar97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 wire694,
                 wire696,
                 (1'h0)};
  assign wire10 = ((!wire8[(1'h0):(1'h0)]) < ($unsigned($signed(wire5)) > $unsigned(wire9[(4'h9):(2'h2)])));
  always
    @(posedge clk) begin
      if (wire6)
        begin
          for (forvar11 = (1'h0); (forvar11 < (2'h2)); forvar11 = (forvar11 + (1'h1)))
            begin
              reg12 <= forvar11[(4'h8):(3'h4)];
            end
          if (wire5)
            begin
              reg13 <= (({wire10[(1'h1):(1'h0)],
                  reg12[(5'h14):(5'h12)]} - $unsigned($signed($signed((8'had))))) ^~ $signed(wire8[(4'h9):(2'h3)]));
              reg14 <= (8'h9c);
            end
          else
            begin
              reg13 <= ((~^$unsigned($signed(((8'hb7) <= reg14)))) >>> wire9);
              reg14 = (8'h9f);
              reg15 <= ($signed("58") ~^ forvar11[(2'h3):(1'h1)]);
            end
          reg16 <= ("ZL0RnD1IAAYd" != (-wire8[(3'h4):(1'h1)]));
          reg17 <= (8'hb1);
          reg18 <= reg14[(4'hd):(4'h8)];
        end
      else
        begin
          for (forvar11 = (1'h0); (forvar11 < (1'h0)); forvar11 = (forvar11 + (1'h1)))
            begin
              reg12 <= reg15[(3'h7):(3'h6)];
              reg13 = {$signed(("nf5797XH4r8NJmon4pB" ?
                      {reg12} : $unsigned((wire7 || (8'ha9))))),
                  {($unsigned(reg12) > (wire5[(1'h1):(1'h0)] >= forvar11))}};
              reg14 <= {reg13};
            end
        end
      for (forvar19 = (1'h0); (forvar19 < (2'h2)); forvar19 = (forvar19 + (1'h1)))
        begin
          for (forvar20 = (1'h0); (forvar20 < (2'h2)); forvar20 = (forvar20 + (1'h1)))
            begin
              reg21 <= forvar19[(3'h6):(3'h4)];
              reg22 <= (8'ha3);
            end
          reg23 = (wire10 ?
              $signed(forvar20[(2'h3):(2'h3)]) : $unsigned($signed((wire10 ~^ $unsigned((8'h9c))))));
        end
      reg24 = reg17[(3'h6):(3'h5)];
      reg25 <= $unsigned({(($unsigned(reg15) || $unsigned(reg17)) != (wire8 ?
              {forvar11} : forvar19[(4'h8):(1'h0)]))});
    end
  always
    @(posedge clk) begin
      if (reg25[(3'h7):(3'h7)])
        begin
          for (forvar26 = (1'h0); (forvar26 < (2'h2)); forvar26 = (forvar26 + (1'h1)))
            begin
              reg27 <= $unsigned($unsigned($unsigned(reg14)));
            end
          reg28 <= (((forvar19[(4'h8):(3'h6)] <<< reg16) ?
              reg21 : (reg27[(4'ha):(3'h7)] ?
                  {wire8,
                      (wire6 || (8'hbf))} : $unsigned(forvar26))) >>> $signed({reg18,
              {(8'hb7), {reg18}}}));
        end
      else
        begin
          reg26 <= (((forvar26[(1'h0):(1'h0)] <= (~^wire8)) ?
              {"h",
                  (8'haf)} : (!forvar11[(1'h0):(1'h0)])) ~^ (~^({$unsigned((8'ha8)),
              ((8'h9f) ? (8'hab) : reg25)} <<< {(reg15 && wire5)})));
          for (forvar27 = (1'h0); (forvar27 < (1'h0)); forvar27 = (forvar27 + (1'h1)))
            begin
              reg28 <= $unsigned(forvar27);
              reg29 = $unsigned(wire7);
              reg30 <= {$signed((($unsigned(reg27) ?
                      $unsigned(wire10) : (wire5 < reg22)) != $unsigned($signed((8'ha4))))),
                  $unsigned($signed((8'hbb)))};
              reg31 <= $unsigned($signed((&"w")));
            end
          for (forvar32 = (1'h0); (forvar32 < (2'h2)); forvar32 = (forvar32 + (1'h1)))
            begin
              reg33 <= $signed((^~("isxHu69XEOLXk04" ?
                  {$unsigned(wire9), (~forvar19)} : reg17)));
              reg34 = wire9[(3'h4):(2'h3)];
              reg35 = $signed({reg34[(4'hc):(4'ha)]});
              reg36 <= wire9[(1'h0):(1'h0)];
            end
        end
      reg37 = forvar11[(4'hb):(4'h8)];
      if (wire9)
        begin
          reg38 = (reg36 >= ({$unsigned($signed(wire6))} > (((~(8'ha5)) * {reg13}) ?
              (~^(!wire6)) : reg26[(3'h4):(3'h4)])));
          reg39 <= forvar11[(4'ha):(4'h9)];
          reg40 <= $signed((reg33 ?
              {(reg22 ? reg27 : reg12[(5'h12):(4'he)]),
                  (reg18 || ((8'had) ? reg30 : forvar32))} : {((reg14 ?
                      (8'haf) : forvar26) - (-reg34)),
                  wire7[(3'h6):(1'h0)]}));
          reg41 <= (reg27[(3'h5):(2'h2)] ?
              reg34 : $signed(($signed(((8'hbe) || forvar26)) == ($unsigned(reg30) >>> reg15[(4'hc):(3'h6)]))));
          reg42 = $unsigned(((^(!(wire10 ? reg26 : reg37))) ?
              $unsigned((7'h41)) : ((reg14 ?
                  $signed(reg18) : $unsigned((7'h44))) ~^ forvar11)));
        end
      else
        begin
          for (forvar38 = (1'h0); (forvar38 < (2'h2)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 = $unsigned($unsigned(wire9));
              reg40 <= ({reg16,
                  reg13} <<< ($signed($unsigned(reg26)) != ((wire7 ?
                      (8'had) : $unsigned(reg22)) ?
                  reg33[(3'h6):(1'h0)] : $signed((-reg34)))));
              reg41 <= ((reg37[(4'h9):(4'h8)] ?
                  (~|(8'ha5)) : ((+(-reg41)) >= ((reg37 ? reg21 : reg27) ?
                      (reg25 ? reg26 : reg24) : reg29))) + reg36);
            end
          reg42 = reg37[(2'h3):(2'h2)];
        end
      for (forvar43 = (1'h0); (forvar43 < (3'h4)); forvar43 = (forvar43 + (1'h1)))
        begin
          for (forvar44 = (1'h0); (forvar44 < (1'h0)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 <= {reg16[(1'h0):(1'h0)]};
              reg46 <= (8'had);
              reg47 <= ($signed("DysMqAi43K9qMLS") >= ($signed({$unsigned(reg42)}) >>> $unsigned({$unsigned((8'haf))})));
            end
        end
    end
  assign wire48 = reg41[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg49 = "PL6OiZV";
      reg50 <= $unsigned(reg39[(4'h8):(3'h7)]);
    end
  assign wire51 = (!($unsigned($unsigned(reg22[(1'h0):(1'h0)])) && {($unsigned((8'ha6)) && wire9[(1'h1):(1'h0)])}));
  always
    @(posedge clk) begin
      reg52 = ({(8'hbc)} >>> ($unsigned(reg26) != ({(8'hbe),
              ((7'h40) ? wire8 : (8'hb9))} ?
          {reg26, (reg35 & reg49)} : reg22[(1'h1):(1'h0)])));
      for (forvar53 = (1'h0); (forvar53 < (2'h2)); forvar53 = (forvar53 + (1'h1)))
        begin
          if ((~|$unsigned(reg42)))
            begin
              reg54 <= forvar19[(3'h4):(2'h2)];
              reg55 = $signed($unsigned($unsigned((((8'h9f) ?
                  reg15 : reg47) << (reg41 < forvar27)))));
              reg56 = $signed(({$unsigned($unsigned((8'hb2)))} < (-forvar27[(3'h5):(2'h3)])));
              reg57 = {(forvar27 || reg42), reg17};
            end
          else
            begin
              reg54 <= reg24;
              reg55 <= ({"9koeNJIt0VP13ftEU"} >= reg50[(5'h12):(3'h6)]);
              reg56 <= (($unsigned($signed((+wire8))) ?
                  $unsigned(($unsigned((7'h40)) ?
                      wire48[(1'h1):(1'h0)] : {forvar27})) : (((reg34 ?
                      reg40 : reg36) >= reg36[(3'h5):(3'h4)]) > ({(8'haa)} - reg49))) & (~^wire48[(1'h1):(1'h0)]));
            end
        end
      for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
        begin
          reg59 = (reg31 ?
              ((reg45[(3'h5):(3'h5)] ?
                  ((wire5 ?
                      reg26 : forvar38) - $unsigned(reg35)) : reg38) - (^~reg33[(3'h4):(3'h4)])) : (8'hb7));
          reg60 <= (^~"J3K4XbAkAdIRwTlQz");
        end
      reg61 = $signed({(7'h44), $signed({$unsigned((7'h41))})});
    end
  always
    @(posedge clk) begin
      reg62 <= $signed(wire5[(1'h0):(1'h0)]);
      for (forvar63 = (1'h0); (forvar63 < (2'h3)); forvar63 = (forvar63 + (1'h1)))
        begin
          reg64 <= reg35;
        end
      reg65 <= (reg31 > $signed(forvar63[(1'h1):(1'h1)]));
      for (forvar66 = (1'h0); (forvar66 < (2'h3)); forvar66 = (forvar66 + (1'h1)))
        begin
          reg67 <= $signed(($unsigned(wire9) ~^ $unsigned($signed({(8'hb4),
              (8'hb7)}))));
          if ($unsigned(reg21))
            begin
              reg68 = (($unsigned(reg61[(3'h4):(3'h4)]) <<< (wire9[(3'h6):(1'h0)] | $unsigned($signed(reg26)))) ?
                  ($unsigned(reg47) * {(8'hb3)}) : {(wire6[(2'h2):(2'h2)] ?
                          ((reg23 == reg13) ? reg12 : reg27) : ((+forvar63) ?
                              {(8'hb6)} : {reg35})),
                      (reg37[(4'hb):(4'ha)] ?
                          wire48[(3'h5):(2'h3)] : ((8'hb6) ?
                              $unsigned(reg42) : wire6[(1'h1):(1'h0)]))});
            end
          else
            begin
              reg68 <= $unsigned(($unsigned(reg25[(1'h0):(1'h0)]) ?
                  (7'h44) : (reg29 == forvar43)));
              reg69 = $signed($signed((!((~&(8'ha9)) ?
                  (reg49 ^ reg38) : {reg30, reg31}))));
              reg70 <= (reg54 ? "OX" : $unsigned($signed((7'h41))));
            end
          for (forvar71 = (1'h0); (forvar71 < (3'h4)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 = "yhPNx";
              reg73 <= reg39[(3'h6):(3'h4)];
            end
          reg74 = {$unsigned(forvar58[(2'h3):(2'h3)]), (forvar11 <<< reg30)};
          for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
            begin
              reg76 <= $signed(((8'hb4) ?
                  (((^forvar27) ?
                      reg72 : ((8'hbb) ?
                          reg69 : reg56)) || forvar26) : ({(reg15 ?
                              reg59 : (8'hb5))} ?
                      (reg14 ?
                          wire8 : $unsigned((8'hae))) : (reg14[(4'he):(2'h2)] ?
                          $unsigned(forvar26) : reg12[(2'h2):(1'h0)]))));
              reg77 <= $signed({wire6, forvar44});
            end
        end
      reg78 = reg52[(4'h8):(4'h8)];
    end
  assign wire79 = (~|$unsigned((&"CzfZh9xIu3Uuip")));
  always
    @(posedge clk) begin
      for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
        begin
          for (forvar81 = (1'h0); (forvar81 < (3'h4)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 <= $unsigned(reg40[(2'h3):(2'h3)]);
              reg83 <= reg72[(2'h2):(1'h1)];
              reg84 = forvar38;
              reg85 <= {{({reg26} + forvar11)}};
            end
          for (forvar86 = (1'h0); (forvar86 < (1'h0)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 <= reg64;
              reg88 <= reg49[(1'h1):(1'h1)];
            end
        end
      for (forvar89 = (1'h0); (forvar89 < (2'h2)); forvar89 = (forvar89 + (1'h1)))
        begin
          for (forvar90 = (1'h0); (forvar90 < (3'h4)); forvar90 = (forvar90 + (1'h1)))
            begin
              reg91 = (~^(reg14 ? forvar86[(3'h6):(2'h2)] : reg85));
              reg92 <= ({$signed((reg56 ?
                          ((8'hb4) || wire51) : $unsigned(forvar86))),
                      forvar53[(4'h8):(3'h4)]} ?
                  $unsigned((reg65 ?
                      (wire79 != ((8'h9f) < (8'ha1))) : (|{forvar86}))) : (~$signed((!((8'hac) >> (8'ha1))))));
              reg93 <= "fOGrzF";
              reg94 = forvar32;
              reg95 = ((forvar44 < forvar19) == (&{(-reg69),
                  {reg31, (reg52 ? (8'h9f) : (8'hb4))}}));
            end
          reg96 <= reg23[(1'h0):(1'h0)];
          for (forvar97 = (1'h0); (forvar97 < (1'h0)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 <= ($unsigned(forvar19) && $unsigned("VAWUyiVEiA4lBmifwYZS"));
              reg99 = ({$signed({$unsigned(forvar43), forvar27}),
                  $signed((8'ha5))} <= reg24);
              reg100 <= ({$signed((8'hb4))} >= reg27[(2'h3):(1'h0)]);
            end
        end
      reg101 = {reg12[(3'h5):(1'h0)]};
      reg102 = forvar27[(5'h10):(5'h10)];
      reg103 <= wire8;
    end
  module104 modinst695 (.wire108(reg77), .y(wire694), .wire107(reg50), .clk(clk), .wire105(reg82), .wire106(reg102));
  module109 modinst697 (wire696, clk, forvar32, reg87, forvar66, reg74, reg61);
  assign wire698 = reg61[(5'h11):(4'he)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module104  (y, clk, wire105, wire106, wire107, wire108);
  output wire [(32'h25e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire105;
  input wire [(5'h10):(1'h0)] wire106;
  input wire signed [(5'h10):(1'h0)] wire107;
  input wire signed [(5'h12):(1'h0)] wire108;
  reg [(5'h12):(1'h0)] reg693 = (1'h0);
  reg [(4'hb):(1'h0)] reg692 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg691 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg690 = (1'h0);
  reg [(2'h3):(1'h0)] reg689 = (1'h0);
  reg [(2'h2):(1'h0)] forvar688 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg687 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar686 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg685 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg684 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg683 = (1'h0);
  reg [(2'h2):(1'h0)] forvar682 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar681 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg680 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg679 = (1'h0);
  reg [(5'h13):(1'h0)] reg678 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg677 = (1'h0);
  reg [(5'h10):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar675 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg674 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg673 = (1'h0);
  reg [(3'h4):(1'h0)] reg672 = (1'h0);
  reg [(4'h9):(1'h0)] reg671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg670 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar669 = (1'h0);
  reg [(4'h9):(1'h0)] reg668 = (1'h0);
  reg [(4'hd):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar666 = (1'h0);
  reg [(2'h3):(1'h0)] forvar665 = (1'h0);
  wire [(4'he):(1'h0)] wire664;
  wire [(4'hd):(1'h0)] wire663;
  wire [(3'h6):(1'h0)] wire661;
  reg [(5'h13):(1'h0)] reg564 = (1'h0);
  reg [(5'h10):(1'h0)] reg563 = (1'h0);
  reg [(4'ha):(1'h0)] reg562 = (1'h0);
  reg signed [(4'he):(1'h0)] reg561 = (1'h0);
  reg [(5'h10):(1'h0)] reg560 = (1'h0);
  reg [(5'h12):(1'h0)] forvar559 = (1'h0);
  reg [(3'h6):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg557 = (1'h0);
  reg [(4'h8):(1'h0)] reg556 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg555 = (1'h0);
  reg [(5'h15):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar552 = (1'h0);
  reg [(5'h13):(1'h0)] reg551 = (1'h0);
  reg [(5'h10):(1'h0)] forvar550 = (1'h0);
  reg [(2'h2):(1'h0)] reg549 = (1'h0);
  reg [(5'h15):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg546 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar545 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire543;
  wire signed [(4'hc):(1'h0)] wire516;
  wire signed [(3'h4):(1'h0)] wire515;
  wire [(5'h11):(1'h0)] wire268;
  wire signed [(3'h7):(1'h0)] wire513;
  assign y = {reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 forvar688,
                 reg687,
                 forvar686,
                 reg685,
                 reg684,
                 reg683,
                 forvar682,
                 forvar681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 forvar675,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 forvar669,
                 reg668,
                 reg667,
                 forvar666,
                 forvar665,
                 wire664,
                 wire663,
                 wire661,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 forvar559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 forvar552,
                 reg551,
                 forvar550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 forvar545,
                 wire543,
                 wire516,
                 wire515,
                 wire268,
                 wire513,
                 (1'h0)};
  module109 modinst269 (wire268, clk, wire105, wire106, wire107, wire108, (8'hb3));
  module270 modinst514 (.wire271(wire108), .wire273(wire106), .y(wire513), .wire272(wire107), .wire274(wire105), .wire275(wire268), .clk(clk));
  assign wire515 = (wire108[(5'h11):(4'hb)] ? wire107 : wire107);
  assign wire516 = (((wire105[(3'h7):(1'h0)] ? {wire515} : $signed(wire268)) ?
                       {$unsigned({wire268, wire515}),
                           $unsigned((~&wire106))} : $unsigned(wire105[(4'ha):(3'h7)])) > ($unsigned(wire108[(4'hb):(3'h6)]) ?
                       ((^wire106) ?
                           ((~^wire105) >= wire268) : (wire513[(1'h0):(1'h0)] > $signed((8'ha8)))) : {wire107,
                           wire108}));
  module517 modinst544 (.wire521(wire513), .y(wire543), .wire519(wire268), .wire520(wire107), .wire518(wire516), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar545 = (1'h0); (forvar545 < (1'h0)); forvar545 = (forvar545 + (1'h1)))
        begin
          reg546 = wire543;
          reg547 <= ((wire105[(2'h3):(1'h0)] * ((8'haa) != wire107[(4'h8):(2'h2)])) >>> ($unsigned({wire268[(4'he):(4'hc)],
              {wire105}}) || {((|wire543) ?
                  $signed(wire108) : $signed(wire106)),
              reg546}));
          reg548 <= wire515[(1'h0):(1'h0)];
          reg549 = {{$unsigned($unsigned($unsigned(reg547)))}};
        end
      for (forvar550 = (1'h0); (forvar550 < (2'h3)); forvar550 = (forvar550 + (1'h1)))
        begin
          reg551 = wire513[(2'h3):(2'h2)];
          for (forvar552 = (1'h0); (forvar552 < (2'h3)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 = $unsigned((($unsigned(reg547[(2'h2):(1'h0)]) ?
                      wire515[(1'h0):(1'h0)] : (-reg549)) ?
                  (($unsigned(wire107) ?
                      (wire515 ~^ (8'ha2)) : $unsigned(wire513)) & $unsigned(reg549)) : (8'hba)));
              reg554 <= ($unsigned((~^$signed((&wire513)))) == wire106[(3'h5):(1'h0)]);
              reg555 <= $unsigned(($unsigned(wire268[(4'hb):(2'h2)]) ?
                  wire516 : wire513));
              reg556 <= $signed((8'ha7));
              reg557 = wire268;
            end
          reg558 = $signed({(($signed((8'ha5)) ?
                  wire515[(1'h0):(1'h0)] : $signed(wire513)) < ((reg554 ?
                  wire106 : (8'ha0)) ^~ reg553[(2'h3):(2'h3)]))});
        end
      for (forvar559 = (1'h0); (forvar559 < (1'h0)); forvar559 = (forvar559 + (1'h1)))
        begin
          reg560 <= $signed($unsigned((|$unsigned($signed(reg557)))));
          reg561 = $unsigned(wire105[(1'h0):(1'h0)]);
          reg562 = (forvar550 <= $unsigned((&reg558[(1'h0):(1'h0)])));
        end
      reg563 <= (^(7'h42));
      reg564 <= wire106;
    end
  module565 modinst662 (wire661, clk, reg557, forvar550, reg563, reg554);
  assign wire663 = (8'hbb);
  assign wire664 = wire516;
  always
    @(posedge clk) begin
      for (forvar665 = (1'h0); (forvar665 < (2'h2)); forvar665 = (forvar665 + (1'h1)))
        begin
          for (forvar666 = (1'h0); (forvar666 < (2'h2)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 <= {(reg555[(2'h2):(1'h1)] ?
                      wire268 : ("M77" & $unsigned($unsigned(wire107))))};
              reg668 <= $signed($unsigned(reg560));
            end
          for (forvar669 = (1'h0); (forvar669 < (1'h0)); forvar669 = (forvar669 + (1'h1)))
            begin
              reg670 <= ((!$unsigned(reg551[(2'h3):(2'h2)])) ?
                  $signed(((~$signed(reg563)) ~^ {(reg668 <<< forvar666)})) : reg557);
              reg671 <= forvar545[(1'h0):(1'h0)];
              reg672 <= (~^(8'ha4));
              reg673 <= (^wire543[(4'hc):(2'h3)]);
              reg674 <= (((wire663 << reg551) >>> (7'h40)) ?
                  wire108[(4'h8):(1'h1)] : reg562[(1'h1):(1'h1)]);
            end
          for (forvar675 = (1'h0); (forvar675 < (3'h4)); forvar675 = (forvar675 + (1'h1)))
            begin
              reg676 <= $unsigned(($signed({forvar552,
                  ((8'hb8) ?
                      reg557 : forvar669)}) & ({reg554[(5'h15):(5'h11)]} && ($unsigned(reg564) - wire105))));
              reg677 = (forvar669[(1'h1):(1'h0)] - $unsigned((!"Dd9")));
              reg678 = reg557;
              reg679 <= ((~&(($unsigned((8'ha2)) ^~ wire513) - wire268)) == $unsigned(forvar665));
              reg680 = ((wire108[(4'h9):(4'h8)] | ((reg668 ?
                  {(8'haf),
                      (7'h40)} : $unsigned(reg561)) >>> {$unsigned(reg671),
                  reg668})) ^ (reg560 >> forvar669));
            end
        end
      for (forvar681 = (1'h0); (forvar681 < (2'h2)); forvar681 = (forvar681 + (1'h1)))
        begin
          for (forvar682 = (1'h0); (forvar682 < (2'h3)); forvar682 = (forvar682 + (1'h1)))
            begin
              reg683 <= wire513[(3'h7):(1'h0)];
            end
          reg684 = wire661;
          reg685 <= $signed({$unsigned($unsigned({wire106, reg547}))});
          for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
            begin
              reg687 <= $unsigned(forvar675[(4'hb):(4'ha)]);
            end
          for (forvar688 = (1'h0); (forvar688 < (1'h1)); forvar688 = (forvar688 + (1'h1)))
            begin
              reg689 <= {{$unsigned($signed({wire515}))},
                  reg667[(3'h6):(3'h5)]};
              reg690 <= forvar545;
              reg691 <= ((+wire515[(1'h0):(1'h0)]) ^~ reg547);
              reg692 = wire664[(4'hb):(3'h4)];
              reg693 = (((8'ha2) ?
                  wire661[(3'h4):(1'h0)] : (^((^~reg549) >>> "G464JtmV"))) + $unsigned(reg673));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module565
#( parameter param660 = ((+{(((8'hb8) ? (8'h9f) : (7'h41)) != ((8'ha9) == (8'hbf))), (|(^(8'haa)))}) ? (((((8'h9d) | (8'ha8)) != {(7'h43)}) ^ ((8'ha3) ? (&(8'hab)) : {(8'hb6), (7'h42)})) + ((7'h43) << (((8'had) << (8'hb5)) < (8'ha9)))) : ((((8'hb5) != ((8'hbd) >= (8'ha5))) >= (&((8'hb6) >>> (8'ha9)))) + (({(8'ha4), (8'ha0)} && (^(8'hb5))) && (((8'hbd) ? (8'haa) : (8'hbf)) ? ((8'hb2) >>> (8'hbb)) : {(8'hba), (8'hb3)})))) )
(y, clk, wire569, wire568, wire567, wire566);
  output wire [(32'h43f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire569;
  input wire [(4'hf):(1'h0)] wire568;
  input wire signed [(4'he):(1'h0)] wire567;
  input wire [(3'h7):(1'h0)] wire566;
  wire signed [(4'hb):(1'h0)] wire659;
  reg [(3'h4):(1'h0)] reg658 = (1'h0);
  reg [(5'h10):(1'h0)] reg657 = (1'h0);
  reg [(5'h12):(1'h0)] reg656 = (1'h0);
  reg [(4'hb):(1'h0)] reg655 = (1'h0);
  reg [(2'h2):(1'h0)] reg654 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg653 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg652 = (1'h0);
  reg [(5'h10):(1'h0)] forvar651 = (1'h0);
  reg [(4'ha):(1'h0)] reg650 = (1'h0);
  reg [(3'h5):(1'h0)] forvar649 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg648 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg647 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire646;
  reg signed [(2'h3):(1'h0)] reg645 = (1'h0);
  reg [(4'h9):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar643 = (1'h0);
  reg [(5'h14):(1'h0)] reg642 = (1'h0);
  reg [(5'h11):(1'h0)] reg641 = (1'h0);
  reg [(5'h11):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg639 = (1'h0);
  reg [(3'h7):(1'h0)] reg638 = (1'h0);
  reg [(3'h7):(1'h0)] reg637 = (1'h0);
  reg [(5'h12):(1'h0)] reg636 = (1'h0);
  reg [(3'h7):(1'h0)] forvar635 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg634 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar633 = (1'h0);
  reg [(4'hc):(1'h0)] reg632 = (1'h0);
  wire signed [(4'he):(1'h0)] wire631;
  wire signed [(4'ha):(1'h0)] wire630;
  wire [(2'h2):(1'h0)] wire629;
  reg signed [(5'h13):(1'h0)] reg628 = (1'h0);
  reg [(4'h9):(1'h0)] reg627 = (1'h0);
  reg [(5'h12):(1'h0)] forvar626 = (1'h0);
  reg [(3'h4):(1'h0)] reg625 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar624 = (1'h0);
  reg [(5'h12):(1'h0)] reg623 = (1'h0);
  reg [(4'hb):(1'h0)] reg622 = (1'h0);
  reg signed [(4'he):(1'h0)] reg621 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar620 = (1'h0);
  reg [(4'ha):(1'h0)] reg619 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar618 = (1'h0);
  reg [(3'h6):(1'h0)] reg617 = (1'h0);
  reg [(3'h4):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg615 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg609 = (1'h0);
  reg [(4'ha):(1'h0)] reg608 = (1'h0);
  reg [(4'hd):(1'h0)] reg607 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg606 = (1'h0);
  reg [(4'h9):(1'h0)] reg605 = (1'h0);
  reg [(3'h4):(1'h0)] reg604 = (1'h0);
  reg [(5'h15):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg602 = (1'h0);
  reg [(5'h10):(1'h0)] reg601 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg600 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg599 = (1'h0);
  reg [(4'ha):(1'h0)] reg598 = (1'h0);
  reg [(4'hd):(1'h0)] reg597 = (1'h0);
  reg [(5'h10):(1'h0)] reg596 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg595 = (1'h0);
  reg [(4'h8):(1'h0)] reg594 = (1'h0);
  reg [(4'hf):(1'h0)] reg593 = (1'h0);
  reg [(3'h4):(1'h0)] reg592 = (1'h0);
  reg [(5'h15):(1'h0)] reg591 = (1'h0);
  reg [(3'h6):(1'h0)] reg590 = (1'h0);
  reg [(4'hb):(1'h0)] forvar589 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar588 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire587;
  reg [(4'h8):(1'h0)] reg586 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg585 = (1'h0);
  reg [(4'h8):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg583 = (1'h0);
  reg [(4'hf):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar580 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg580 = (1'h0);
  wire [(2'h3):(1'h0)] wire579;
  wire signed [(3'h5):(1'h0)] wire578;
  wire signed [(5'h13):(1'h0)] wire577;
  wire [(4'ha):(1'h0)] wire576;
  wire [(5'h10):(1'h0)] wire575;
  wire signed [(4'hd):(1'h0)] wire574;
  wire signed [(4'hf):(1'h0)] wire573;
  wire [(5'h11):(1'h0)] wire572;
  wire signed [(3'h6):(1'h0)] wire571;
  wire signed [(5'h12):(1'h0)] wire570;
  assign y = {wire659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 forvar651,
                 reg650,
                 forvar649,
                 reg648,
                 reg647,
                 wire646,
                 reg645,
                 reg644,
                 forvar643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 forvar635,
                 reg634,
                 forvar633,
                 reg632,
                 wire631,
                 wire630,
                 wire629,
                 reg628,
                 reg627,
                 forvar626,
                 reg625,
                 forvar624,
                 reg623,
                 reg622,
                 reg621,
                 forvar620,
                 reg619,
                 forvar618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 forvar589,
                 forvar588,
                 wire587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 forvar580,
                 reg580,
                 wire579,
                 wire578,
                 wire577,
                 wire576,
                 wire575,
                 wire574,
                 wire573,
                 wire572,
                 wire571,
                 wire570,
                 (1'h0)};
  assign wire570 = wire567;
  assign wire571 = wire567;
  assign wire572 = (wire568[(3'h6):(1'h1)] - (wire569 ^~ wire571[(2'h2):(1'h1)]));
  assign wire573 = $unsigned((8'h9d));
  assign wire574 = wire569;
  assign wire575 = (^~$unsigned($unsigned($unsigned(wire566))));
  assign wire576 = ((8'ha6) > (wire575 & $signed({(|(8'ha8))})));
  assign wire577 = (($unsigned($signed(wire576[(3'h5):(1'h1)])) ~^ ((wire571[(3'h4):(1'h0)] <= $unsigned(wire575)) << wire576)) || ({wire574} <<< (wire571 ?
                       {(wire574 & wire571)} : $unsigned((wire571 < wire569)))));
  assign wire578 = wire575;
  assign wire579 = "Pgud9dMz";
  always
    @(posedge clk) begin
      if ((wire578[(3'h5):(3'h4)] >> ((($unsigned(wire578) ^~ wire566[(3'h7):(2'h3)]) * (wire579 ?
              wire568 : wire570[(2'h3):(1'h0)])) ?
          (wire573 ? wire568[(4'he):(4'ha)] : wire569) : wire577)))
        begin
          reg580 <= wire566[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar580 = (1'h0); (forvar580 < (3'h4)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg581 = (8'hb8);
            end
          reg582 <= {wire574, wire570};
          reg583 <= reg580;
        end
      reg584 <= (~|forvar580);
      reg585 = (8'hbd);
      reg586 <= (({wire573,
          ({reg585} - {(8'ha8)})} && (8'h9f)) & $unsigned(({reg584[(3'h4):(3'h4)],
          (wire573 & wire566)} + {wire572, {(8'ha2), wire567}})));
    end
  assign wire587 = {{wire571}};
  always
    @(posedge clk) begin
      for (forvar588 = (1'h0); (forvar588 < (3'h4)); forvar588 = (forvar588 + (1'h1)))
        begin
          for (forvar589 = (1'h0); (forvar589 < (2'h2)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 <= ($signed($unsigned((((8'hb0) || wire574) & $signed((8'hb1))))) >= (({(~|wire569)} > $unsigned(wire571)) ?
                  ($unsigned((reg585 ?
                      wire571 : wire573)) <<< forvar589[(3'h4):(2'h2)]) : (^wire570[(4'hf):(4'h9)])));
              reg591 = $unsigned((8'had));
              reg592 = (~^reg591);
              reg593 = {(8'hbf)};
              reg594 = (8'haf);
            end
        end
      reg595 = ($signed($unsigned(reg590[(3'h5):(1'h0)])) ?
          ({{forvar589[(1'h1):(1'h0)], $signed((8'ha1))}} ?
              ($unsigned($signed(reg586)) || $signed((wire574 == reg585))) : (8'ha6)) : ((7'h42) < $unsigned(wire572)));
      if ({((((reg586 ^ reg592) >= ((8'h9e) ? (8'hb5) : wire567)) & {reg593,
              reg591[(5'h10):(3'h5)]}) << $unsigned(wire571[(1'h0):(1'h0)]))})
        begin
          if ($unsigned(wire571[(3'h5):(3'h4)]))
            begin
              reg596 <= ($unsigned({(!wire578)}) ? wire579 : reg594);
              reg597 <= {(forvar588 ?
                      wire575[(4'ha):(2'h3)] : ($signed((^wire574)) ?
                          forvar589 : wire574)),
                  reg581[(3'h7):(2'h3)]};
              reg598 <= (~^((reg580[(4'hc):(2'h2)] <<< (7'h44)) ?
                  $unsigned({$unsigned((8'had)),
                      (~&forvar588)}) : $unsigned($unsigned((reg583 ^ (8'hb3))))));
              reg599 = reg597;
            end
          else
            begin
              reg596 = $unsigned($signed(reg599));
            end
          reg600 = $signed((8'hbc));
        end
      else
        begin
          reg596 <= {(-wire577[(4'ha):(3'h4)])};
        end
      reg601 <= (((7'h44) ?
              ((reg596[(4'ha):(4'h9)] && {(8'hba),
                  forvar580}) >= wire568) : reg580[(3'h5):(1'h1)]) ?
          (&(reg596[(4'hd):(4'ha)] ?
              {reg596[(5'h10):(4'ha)]} : {reg595[(3'h5):(1'h0)],
                  $unsigned((8'h9d))})) : wire579);
      if (forvar580)
        begin
          reg602 <= wire587;
          reg603 = $signed(((~&{(wire578 | (8'hbc))}) ?
              {$signed((reg581 < wire575)),
                  ($signed((8'hb9)) ?
                      reg591[(1'h1):(1'h0)] : $unsigned(reg594))} : {reg592,
                  $unsigned(((8'ha4) ? (8'hb7) : reg590))}));
        end
      else
        begin
          if (((((&reg584) ?
              ((8'ha1) + (wire566 <<< (8'haf))) : {((8'hb6) >= reg592),
                  {(8'ha0)}}) ^~ {wire577, {(wire577 >>> reg582)}}) < reg602))
            begin
              reg602 = {forvar588[(4'hb):(3'h4)]};
            end
          else
            begin
              reg602 <= (({(reg594 != wire575[(3'h5):(2'h3)]),
                  forvar589[(4'hb):(4'ha)]} != (~&((reg586 <= reg590) >>> {(7'h42)}))) >>> {$unsigned((wire577 | forvar580))});
              reg603 = ({($signed($signed(reg601)) ?
                          (reg583 ?
                              (reg596 ?
                                  reg594 : reg580) : (reg590 > wire579)) : {reg583,
                              reg586[(1'h1):(1'h1)]})} ?
                  {((~^$unsigned((8'hba))) < $unsigned($unsigned((8'hb7))))} : ({wire575} ?
                      reg601 : "CSfsYCXp2u908C"));
              reg604 = $unsigned({reg583, reg593});
              reg605 = $unsigned($unsigned(reg602[(4'h8):(3'h5)]));
            end
          reg606 = "hpPT6sTRHeuC";
          reg607 <= (8'ha5);
          if ($unsigned(($unsigned($signed((reg591 ?
              (8'had) : (7'h42)))) ^~ reg580[(5'h11):(4'hd)])))
            begin
              reg608 <= $unsigned(wire571[(2'h2):(1'h1)]);
              reg609 <= $unsigned(reg606[(4'hd):(2'h2)]);
              reg610 <= ($unsigned((^~$unsigned((8'ha1)))) ?
                  {(8'hb1)} : $unsigned((8'h9c)));
            end
          else
            begin
              reg608 <= reg585;
              reg609 = $unsigned($unsigned(reg593[(3'h5):(2'h2)]));
              reg610 = reg599;
              reg611 <= {(8'hb2)};
              reg612 <= {(8'hb6),
                  $unsigned($signed({$signed(wire576), "D2G1fmQMeI"}))};
            end
        end
    end
  always
    @(posedge clk) begin
      reg613 <= wire569;
      reg614 <= reg591;
      reg615 = (reg599[(3'h4):(1'h0)] - reg600[(1'h0):(1'h0)]);
      reg616 <= (reg580 ^ (8'ha6));
    end
  always
    @(posedge clk) begin
      reg617 <= wire578;
      for (forvar618 = (1'h0); (forvar618 < (2'h3)); forvar618 = (forvar618 + (1'h1)))
        begin
          reg619 <= $unsigned(($unsigned((reg594 ? reg593 : (~&wire566))) ?
              (~reg609[(4'hd):(1'h0)]) : wire566[(1'h0):(1'h0)]));
        end
      for (forvar620 = (1'h0); (forvar620 < (3'h4)); forvar620 = (forvar620 + (1'h1)))
        begin
          reg621 = {$unsigned((8'h9e)), forvar618};
          reg622 = reg581;
        end
      reg623 <= reg585;
      for (forvar624 = (1'h0); (forvar624 < (1'h1)); forvar624 = (forvar624 + (1'h1)))
        begin
          reg625 = reg619[(4'h9):(4'h9)];
          for (forvar626 = (1'h0); (forvar626 < (1'h0)); forvar626 = (forvar626 + (1'h1)))
            begin
              reg627 <= $unsigned({"nRX5CfWi"});
              reg628 <= (8'ha4);
            end
        end
    end
  assign wire629 = reg582;
  assign wire630 = forvar626;
  assign wire631 = reg590[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg632 <= ((~|reg594[(4'h8):(3'h4)]) == "5IC");
      for (forvar633 = (1'h0); (forvar633 < (1'h0)); forvar633 = (forvar633 + (1'h1)))
        begin
          reg634 <= $signed($unsigned((reg622[(4'h9):(3'h6)] | {$signed(wire570),
              $unsigned((8'hb4))})));
          for (forvar635 = (1'h0); (forvar635 < (2'h2)); forvar635 = (forvar635 + (1'h1)))
            begin
              reg636 = (({((wire574 & reg590) || wire568[(4'hb):(2'h3)]),
                      wire576} || {(8'hb2), $unsigned($unsigned(wire568))}) ?
                  wire577[(5'h10):(4'h8)] : wire630);
              reg637 = reg593[(2'h3):(2'h3)];
              reg638 = reg625;
            end
          reg639 <= (((8'ha3) >> "U9Iud7g3xkr6W1") ?
              ($unsigned(((8'hbd) * {wire567,
                  reg582})) >= $signed({reg610[(3'h6):(3'h6)]})) : ($unsigned(($signed(reg605) <<< ((8'hb4) && forvar635))) ?
                  (&reg602[(2'h3):(2'h2)]) : $unsigned(({reg591} ?
                      wire567 : $unsigned(reg586)))));
          reg640 <= reg600;
          if (forvar620[(4'hd):(4'h9)])
            begin
              reg641 = (8'hbf);
            end
          else
            begin
              reg641 <= $signed($unsigned($signed(forvar633[(4'ha):(4'h9)])));
              reg642 <= ((~^reg614[(4'hd):(3'h6)]) - ((!"ZbiORYgPDm7NmCbT") > {({(8'h9e),
                      forvar588} | "")}));
            end
        end
      for (forvar643 = (1'h0); (forvar643 < (2'h3)); forvar643 = (forvar643 + (1'h1)))
        begin
          reg644 = reg612[(4'h8):(1'h1)];
          reg645 = {{{reg622[(2'h3):(2'h2)]}, reg592[(1'h0):(1'h0)]}, (8'ha4)};
        end
    end
  assign wire646 = $unsigned($signed({{{forvar620, wire576}}, reg599}));
  always
    @(posedge clk) begin
      reg647 = ((reg585[(2'h3):(1'h1)] <= $signed(($signed(reg596) ^ $unsigned((8'hac))))) ?
          ({wire587[(3'h4):(2'h2)],
              wire629} < (&{(reg614 ~^ forvar618)})) : (8'hb4));
      reg648 <= ($unsigned($unsigned((~|forvar624))) > (~|$unsigned(reg636[(4'hf):(1'h0)])));
      for (forvar649 = (1'h0); (forvar649 < (1'h1)); forvar649 = (forvar649 + (1'h1)))
        begin
          reg650 = reg593;
          for (forvar651 = (1'h0); (forvar651 < (2'h3)); forvar651 = (forvar651 + (1'h1)))
            begin
              reg652 <= {((forvar620[(3'h4):(2'h2)] - $unsigned($unsigned(reg615))) ?
                      (wire569 ?
                          (wire576 << $unsigned((8'haa))) : ((wire578 ?
                              wire572 : forvar635) < (forvar643 ?
                              (7'h44) : reg590))) : $signed(reg595[(1'h0):(1'h0)])),
                  (wire579[(2'h3):(2'h3)] <= reg606)};
              reg653 <= $unsigned($unsigned($unsigned($signed(((8'h9f) <<< (8'hbd))))));
              reg654 <= $signed(reg603);
              reg655 <= (((8'hbb) ?
                  reg619[(3'h5):(1'h0)] : $unsigned((8'ha5))) ^~ $unsigned((^(7'h43))));
              reg656 = (reg595 + (^{(wire630[(4'ha):(4'ha)] <= (-(8'ha2))),
                  (reg605[(3'h4):(2'h3)] ?
                      ((8'ha1) >= reg632) : $unsigned(reg606))}));
            end
        end
      reg657 <= $unsigned((7'h44));
      reg658 <= {"b6MNuhf"};
    end
  assign wire659 = reg650[(2'h2):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module517
#( parameter param541 = ((((~&((8'haf) | (8'h9f))) < (((8'hab) ? (8'ha7) : (7'h41)) >= ((7'h40) ? (8'hb4) : (8'ha8)))) <<< ((((8'hbe) ? (8'haa) : (7'h43)) & ((8'h9d) <<< (7'h44))) ? (-((8'ha4) >> (8'hb0))) : ({(8'hbe), (8'hb8)} ? {(8'hb9)} : ((8'hab) ? (8'hb0) : (8'ha2))))) ? ((&(-((8'had) ? (8'ha5) : (8'hbc)))) * (&(&{(8'ha9), (8'hba)}))) : ((+(7'h44)) & {(8'hb0)}))
, parameter param542 = ((|(((param541 >= param541) << (param541 == param541)) ? param541 : {param541, (param541 ? param541 : param541)})) ? (~(param541 && param541)) : (+(({param541} > (~|(8'ha5))) ? {(+(8'hb1)), (param541 <= (8'hac))} : (((8'hb2) ? (8'hbb) : param541) > ((8'h9f) ? param541 : (7'h42)))))) )
(y, clk, wire521, wire520, wire519, wire518);
  output wire [(32'hee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire521;
  input wire signed [(5'h10):(1'h0)] wire520;
  input wire [(4'he):(1'h0)] wire519;
  input wire signed [(4'hb):(1'h0)] wire518;
  wire [(5'h11):(1'h0)] wire540;
  wire signed [(2'h2):(1'h0)] wire539;
  wire [(5'h11):(1'h0)] wire538;
  wire signed [(5'h12):(1'h0)] wire537;
  reg signed [(3'h4):(1'h0)] reg536 = (1'h0);
  wire [(4'hc):(1'h0)] wire535;
  wire [(5'h15):(1'h0)] wire534;
  reg signed [(5'h10):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg531 = (1'h0);
  reg [(2'h2):(1'h0)] reg530 = (1'h0);
  reg [(3'h7):(1'h0)] reg529 = (1'h0);
  reg [(4'hd):(1'h0)] reg528 = (1'h0);
  reg [(4'hf):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg526 = (1'h0);
  reg [(3'h7):(1'h0)] reg525 = (1'h0);
  reg [(5'h14):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar523 = (1'h0);
  reg [(5'h10):(1'h0)] reg522 = (1'h0);
  assign y = {wire540,
                 wire539,
                 wire538,
                 wire537,
                 reg536,
                 wire535,
                 wire534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 forvar523,
                 reg522,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg522 = wire521;
    end
  always
    @(posedge clk) begin
      for (forvar523 = (1'h0); (forvar523 < (3'h4)); forvar523 = (forvar523 + (1'h1)))
        begin
          if ((((wire519[(3'h4):(3'h4)] ?
              ($signed(reg522) ^ $signed(reg522)) : (wire519[(3'h6):(3'h5)] <<< (wire521 ?
                  wire520 : wire519))) & $unsigned((((8'haf) && wire520) ~^ forvar523[(5'h14):(4'hc)]))) >>> ((wire518[(4'h9):(3'h4)] << $unsigned(wire519)) ?
              (reg522[(1'h1):(1'h0)] >>> wire518[(3'h6):(1'h0)]) : ({(8'haf)} ?
                  (&$unsigned((8'had))) : $unsigned({forvar523, (8'ha7)})))))
            begin
              reg524 <= {{reg522},
                  (((-(^(8'hb3))) <<< wire520) ?
                      wire518 : ($unsigned((wire519 || forvar523)) | wire518))};
              reg525 = wire520[(4'hf):(3'h5)];
              reg526 = "zZlur0Z5quXGn";
              reg527 <= wire518[(3'h7):(1'h1)];
              reg528 <= $unsigned(wire519);
            end
          else
            begin
              reg524 <= wire519[(2'h2):(2'h2)];
              reg525 <= {(({(&reg528)} + wire521[(2'h3):(2'h3)]) < reg527)};
              reg526 = reg526;
              reg527 <= ((((&((8'hb0) ^ reg522)) << {((8'ha7) <= reg527)}) <= reg527[(1'h1):(1'h1)]) >>> {forvar523,
                  (wire519 > $unsigned(((8'hb5) != wire518)))});
            end
          reg529 <= wire521;
          reg530 <= (((^~$unsigned(reg527)) < (wire518[(3'h4):(3'h4)] ~^ $unsigned((8'hba)))) <<< (8'had));
          reg531 <= reg527[(3'h6):(2'h3)];
        end
      reg532 <= ($unsigned($signed(((reg529 || reg522) >>> (8'h9d)))) >>> reg526[(3'h5):(1'h0)]);
      reg533 <= (~(reg528[(3'h4):(2'h2)] <<< (~&{reg526, (~reg532)})));
    end
  assign wire534 = reg530[(1'h1):(1'h1)];
  assign wire535 = $signed(wire518[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      reg536 <= {reg527[(4'h9):(3'h6)]};
    end
  assign wire537 = (((((7'h44) <<< {(8'ha8)}) ?
                               $unsigned(((8'ha7) ?
                                   wire518 : wire520)) : ("IykL" ?
                                   wire534 : (reg525 >>> (8'hb9)))) ?
                           (-(reg532[(3'h6):(3'h5)] >= reg526)) : wire519) ?
                       (($signed(reg522) <= reg528[(1'h0):(1'h0)]) != (8'had)) : wire520);
  assign wire538 = reg524[(4'hd):(3'h6)];
  assign wire539 = (($unsigned((-reg530)) ?
                       $unsigned($unsigned($signed(reg526))) : wire521) & forvar523[(5'h14):(4'he)]);
  assign wire540 = (wire520 ?
                       $signed(wire519[(4'hb):(3'h6)]) : (($unsigned((8'hae)) && $signed($signed(reg529))) ~^ (reg525[(2'h3):(2'h2)] || reg536[(1'h0):(1'h0)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module270  (y, clk, wire275, wire274, wire273, wire272, wire271);
  output wire [(32'hb1d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire275;
  input wire [(3'h6):(1'h0)] wire274;
  input wire [(5'h10):(1'h0)] wire273;
  input wire signed [(4'h9):(1'h0)] wire272;
  input wire signed [(4'hb):(1'h0)] wire271;
  wire [(3'h6):(1'h0)] wire512;
  wire [(5'h15):(1'h0)] wire511;
  wire [(5'h11):(1'h0)] wire510;
  reg signed [(4'hf):(1'h0)] reg509 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg508 = (1'h0);
  reg [(3'h6):(1'h0)] reg507 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar506 = (1'h0);
  reg [(3'h4):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg504 = (1'h0);
  reg [(3'h7):(1'h0)] forvar503 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg502 = (1'h0);
  reg [(4'hd):(1'h0)] reg501 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg500 = (1'h0);
  reg [(5'h11):(1'h0)] reg499 = (1'h0);
  reg [(5'h15):(1'h0)] forvar498 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg497 = (1'h0);
  reg [(5'h14):(1'h0)] reg496 = (1'h0);
  reg [(5'h12):(1'h0)] forvar495 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg494 = (1'h0);
  reg [(5'h14):(1'h0)] reg493 = (1'h0);
  reg [(4'hc):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg491 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg490 = (1'h0);
  reg [(4'h9):(1'h0)] reg489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg488 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg487 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar486 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg485 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg484 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg483 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg481 = (1'h0);
  reg [(5'h11):(1'h0)] forvar480 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg478 = (1'h0);
  reg [(4'hc):(1'h0)] reg477 = (1'h0);
  reg [(2'h3):(1'h0)] reg476 = (1'h0);
  wire [(3'h6):(1'h0)] wire475;
  reg [(4'hf):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg473 = (1'h0);
  reg [(2'h3):(1'h0)] reg472 = (1'h0);
  reg [(5'h11):(1'h0)] reg471 = (1'h0);
  reg [(4'ha):(1'h0)] forvar470 = (1'h0);
  reg [(4'hd):(1'h0)] reg469 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg468 = (1'h0);
  reg [(5'h13):(1'h0)] reg467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg466 = (1'h0);
  reg [(4'h9):(1'h0)] forvar465 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg464 = (1'h0);
  reg [(4'h8):(1'h0)] reg463 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg462 = (1'h0);
  reg [(3'h5):(1'h0)] reg461 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg460 = (1'h0);
  reg [(4'h8):(1'h0)] forvar459 = (1'h0);
  reg [(5'h13):(1'h0)] reg458 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg457 = (1'h0);
  reg [(3'h6):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar455 = (1'h0);
  reg [(4'hf):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg453 = (1'h0);
  reg [(3'h7):(1'h0)] forvar452 = (1'h0);
  wire [(5'h14):(1'h0)] wire451;
  wire [(2'h2):(1'h0)] wire450;
  reg [(5'h15):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg444 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg448 = (1'h0);
  reg [(2'h3):(1'h0)] reg447 = (1'h0);
  reg [(2'h2):(1'h0)] reg446 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg445 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar444 = (1'h0);
  reg [(4'he):(1'h0)] reg443 = (1'h0);
  reg [(5'h12):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg441 = (1'h0);
  reg [(4'ha):(1'h0)] reg440 = (1'h0);
  reg [(5'h12):(1'h0)] reg439 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg438 = (1'h0);
  reg [(4'ha):(1'h0)] reg437 = (1'h0);
  reg [(4'he):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg435 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg434 = (1'h0);
  reg [(5'h14):(1'h0)] reg433 = (1'h0);
  reg [(5'h13):(1'h0)] reg432 = (1'h0);
  reg [(5'h15):(1'h0)] forvar431 = (1'h0);
  reg [(2'h3):(1'h0)] reg430 = (1'h0);
  reg [(4'hb):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg428 = (1'h0);
  reg [(5'h10):(1'h0)] reg427 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg426 = (1'h0);
  reg [(4'hc):(1'h0)] forvar425 = (1'h0);
  reg signed [(4'he):(1'h0)] reg424 = (1'h0);
  reg [(4'hd):(1'h0)] reg423 = (1'h0);
  reg [(3'h6):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg420 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar419 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar418 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg417 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg415 = (1'h0);
  reg [(4'h9):(1'h0)] reg414 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg407 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar405 = (1'h0);
  reg [(4'h8):(1'h0)] reg403 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg412 = (1'h0);
  reg [(4'ha):(1'h0)] reg411 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg410 = (1'h0);
  reg [(4'h9):(1'h0)] reg409 = (1'h0);
  reg [(3'h7):(1'h0)] reg408 = (1'h0);
  reg [(3'h6):(1'h0)] forvar407 = (1'h0);
  reg [(3'h4):(1'h0)] reg406 = (1'h0);
  reg [(5'h12):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg404 = (1'h0);
  reg [(5'h13):(1'h0)] forvar403 = (1'h0);
  reg [(5'h15):(1'h0)] forvar388 = (1'h0);
  reg [(4'hb):(1'h0)] reg402 = (1'h0);
  reg [(2'h3):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg400 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg398 = (1'h0);
  reg [(5'h15):(1'h0)] reg397 = (1'h0);
  reg [(2'h2):(1'h0)] reg396 = (1'h0);
  reg [(4'hc):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg394 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar393 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg392 = (1'h0);
  reg [(4'h8):(1'h0)] reg391 = (1'h0);
  reg [(5'h10):(1'h0)] reg390 = (1'h0);
  reg [(5'h14):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg388 = (1'h0);
  reg [(4'hb):(1'h0)] reg387 = (1'h0);
  wire [(5'h14):(1'h0)] wire386;
  wire [(4'hb):(1'h0)] wire385;
  wire signed [(5'h10):(1'h0)] wire384;
  reg signed [(2'h2):(1'h0)] reg383 = (1'h0);
  reg [(4'hc):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg370 = (1'h0);
  reg signed [(4'he):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg380 = (1'h0);
  reg [(2'h2):(1'h0)] reg379 = (1'h0);
  reg [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg376 = (1'h0);
  reg [(2'h3):(1'h0)] reg375 = (1'h0);
  reg [(5'h11):(1'h0)] reg374 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg373 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar372 = (1'h0);
  reg [(2'h3):(1'h0)] reg371 = (1'h0);
  reg [(4'h9):(1'h0)] forvar370 = (1'h0);
  reg [(3'h5):(1'h0)] reg369 = (1'h0);
  reg signed [(4'he):(1'h0)] reg368 = (1'h0);
  reg [(4'hc):(1'h0)] reg367 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar366 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar365 = (1'h0);
  reg [(4'h9):(1'h0)] reg364 = (1'h0);
  reg [(3'h7):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg362 = (1'h0);
  reg [(5'h13):(1'h0)] reg361 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg360 = (1'h0);
  reg [(3'h6):(1'h0)] reg359 = (1'h0);
  reg [(5'h13):(1'h0)] reg358 = (1'h0);
  reg [(4'ha):(1'h0)] forvar357 = (1'h0);
  reg [(5'h10):(1'h0)] reg352 = (1'h0);
  reg [(5'h13):(1'h0)] forvar351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg356 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg355 = (1'h0);
  reg [(4'he):(1'h0)] reg354 = (1'h0);
  reg [(4'hc):(1'h0)] reg353 = (1'h0);
  reg [(4'h9):(1'h0)] forvar352 = (1'h0);
  reg [(5'h14):(1'h0)] reg351 = (1'h0);
  reg [(4'h9):(1'h0)] reg350 = (1'h0);
  reg signed [(4'he):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg348 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg347 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg346 = (1'h0);
  reg [(2'h2):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg344 = (1'h0);
  reg [(5'h10):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar342 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg341 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar340 = (1'h0);
  reg [(3'h6):(1'h0)] reg339 = (1'h0);
  reg [(2'h2):(1'h0)] reg338 = (1'h0);
  reg [(4'he):(1'h0)] reg337 = (1'h0);
  reg [(4'hc):(1'h0)] reg336 = (1'h0);
  reg [(4'hd):(1'h0)] forvar335 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg334 = (1'h0);
  reg [(3'h4):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg332 = (1'h0);
  reg [(5'h13):(1'h0)] forvar331 = (1'h0);
  reg [(5'h12):(1'h0)] reg330 = (1'h0);
  reg [(4'he):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg328 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg327 = (1'h0);
  reg signed [(4'he):(1'h0)] reg326 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg325 = (1'h0);
  reg [(4'ha):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg323 = (1'h0);
  reg [(5'h13):(1'h0)] forvar322 = (1'h0);
  reg [(4'hd):(1'h0)] reg321 = (1'h0);
  reg [(4'h8):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar319 = (1'h0);
  reg [(5'h13):(1'h0)] forvar318 = (1'h0);
  reg [(3'h6):(1'h0)] reg317 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg316 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg314 = (1'h0);
  reg [(3'h7):(1'h0)] reg313 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg312 = (1'h0);
  reg [(5'h14):(1'h0)] reg311 = (1'h0);
  reg [(3'h4):(1'h0)] reg310 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg308 = (1'h0);
  reg [(5'h15):(1'h0)] reg307 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar306 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg305 = (1'h0);
  reg [(4'ha):(1'h0)] forvar304 = (1'h0);
  reg [(5'h10):(1'h0)] reg303 = (1'h0);
  reg [(5'h14):(1'h0)] reg302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg301 = (1'h0);
  reg [(3'h5):(1'h0)] forvar300 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg299 = (1'h0);
  reg [(4'hc):(1'h0)] reg298 = (1'h0);
  reg [(4'hc):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg296 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg295 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg294 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg [(4'he):(1'h0)] forvar292 = (1'h0);
  reg [(4'h8):(1'h0)] reg291 = (1'h0);
  reg [(4'he):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg288 = (1'h0);
  reg [(3'h4):(1'h0)] forvar287 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar279 = (1'h0);
  reg [(4'hb):(1'h0)] reg277 = (1'h0);
  reg [(3'h5):(1'h0)] reg289 = (1'h0);
  reg [(5'h12):(1'h0)] forvar288 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg286 = (1'h0);
  reg [(4'hd):(1'h0)] forvar285 = (1'h0);
  reg [(4'hf):(1'h0)] reg284 = (1'h0);
  reg [(5'h12):(1'h0)] reg283 = (1'h0);
  reg [(4'ha):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg281 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg280 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar277 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire276;
  assign y = {wire512,
                 wire511,
                 wire510,
                 reg509,
                 reg508,
                 reg507,
                 forvar506,
                 reg505,
                 reg504,
                 forvar503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 forvar498,
                 reg497,
                 reg496,
                 forvar495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 forvar486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 wire475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 forvar465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 forvar459,
                 reg458,
                 reg457,
                 reg456,
                 forvar455,
                 reg454,
                 reg453,
                 forvar452,
                 wire451,
                 wire450,
                 reg449,
                 reg444,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 forvar444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 forvar431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 forvar425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 forvar419,
                 forvar418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg407,
                 forvar405,
                 reg403,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 reg405,
                 reg404,
                 forvar403,
                 forvar388,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 wire386,
                 wire385,
                 wire384,
                 reg383,
                 reg372,
                 reg370,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 forvar372,
                 reg371,
                 forvar370,
                 reg369,
                 reg368,
                 reg367,
                 forvar366,
                 forvar365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 forvar357,
                 reg352,
                 forvar351,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 forvar352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 forvar342,
                 reg341,
                 forvar340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 forvar335,
                 reg334,
                 reg333,
                 reg332,
                 forvar331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 forvar322,
                 reg321,
                 reg320,
                 forvar319,
                 forvar318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 forvar306,
                 reg305,
                 forvar304,
                 reg303,
                 reg302,
                 reg301,
                 forvar300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 forvar292,
                 reg291,
                 reg290,
                 reg288,
                 forvar287,
                 forvar279,
                 reg277,
                 reg289,
                 forvar288,
                 reg287,
                 reg286,
                 forvar285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 forvar277,
                 wire276,
                 (1'h0)};
  assign wire276 = wire275;
  always
    @(posedge clk) begin
      if (wire276[(1'h1):(1'h0)])
        begin
          for (forvar277 = (1'h0); (forvar277 < (1'h0)); forvar277 = (forvar277 + (1'h1)))
            begin
              reg278 = {{wire276, (8'haa)},
                  {forvar277[(2'h2):(2'h2)], (8'ha2)}};
              reg279 = $unsigned(wire275[(4'ha):(3'h4)]);
            end
          if (wire274)
            begin
              reg280 <= (|((8'ha2) <<< $unsigned(wire273)));
              reg281 <= wire272;
              reg282 = ((-(~forvar277)) | $signed(forvar277));
              reg283 <= ({((+wire273[(2'h2):(2'h2)]) | ((reg281 <<< reg282) < $unsigned((8'hb2))))} > $unsigned({((8'hb3) ?
                      $signed(wire275) : $signed((7'h42)))}));
              reg284 <= reg283[(4'he):(3'h4)];
            end
          else
            begin
              reg280 <= wire274;
              reg281 <= {$signed(((!(-(8'hb9))) ?
                      $signed(reg283) : (+(reg280 ^~ wire273))))};
              reg282 = $signed((((forvar277 ?
                  reg278[(4'hf):(3'h6)] : reg280[(1'h0):(1'h0)]) >>> reg279[(1'h1):(1'h0)]) & $signed(wire275)));
            end
          for (forvar285 = (1'h0); (forvar285 < (1'h1)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 <= (8'hac);
              reg287 <= ({$signed(wire271[(3'h7):(1'h1)])} ?
                  (($signed(reg282) + (((8'hbd) ^ wire271) ?
                      (wire272 ~^ (8'hab)) : {(8'hb9)})) > (wire271[(2'h2):(1'h0)] ^ (+{reg284,
                      reg279}))) : reg283);
            end
          for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
            begin
              reg289 <= {$unsigned($unsigned("zam"))};
            end
        end
      else
        begin
          reg277 <= $unsigned($unsigned((($unsigned((8'hb5)) ?
                  (~|(7'h40)) : reg282[(3'h6):(1'h0)]) ?
              reg280 : (&(-(8'ha5))))));
          reg278 <= (!($signed($unsigned(((7'h43) ~^ wire273))) ~^ ((8'hb2) | reg278[(2'h2):(1'h1)])));
          for (forvar279 = (1'h0); (forvar279 < (2'h3)); forvar279 = (forvar279 + (1'h1)))
            begin
              reg280 <= $unsigned(forvar277[(1'h1):(1'h0)]);
              reg281 <= wire274[(2'h2):(2'h2)];
              reg282 <= {{{{forvar288}, wire272[(4'h9):(2'h2)]},
                      $signed((7'h41))},
                  ($unsigned(reg289) & $signed(wire272[(4'h9):(3'h5)]))};
              reg283 <= $unsigned({$signed((&(-wire271))),
                  {(|wire275), (reg283 ? wire271[(3'h6):(2'h3)] : {reg277})}});
              reg284 = (8'hb3);
            end
          for (forvar285 = (1'h0); (forvar285 < (2'h3)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 <= (reg278 + (wire272 ?
                  {reg281[(1'h0):(1'h0)]} : forvar288));
            end
          for (forvar287 = (1'h0); (forvar287 < (2'h2)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 <= (8'h9d);
              reg289 <= {(|forvar288)};
              reg290 <= ($unsigned($signed($unsigned(forvar287))) + {{{reg284[(4'h8):(2'h3)]}}});
              reg291 = reg289;
            end
        end
      for (forvar292 = (1'h0); (forvar292 < (1'h1)); forvar292 = (forvar292 + (1'h1)))
        begin
          reg293 <= {reg287};
          reg294 <= $signed("rBZayC96");
          if ($signed(reg284[(4'h9):(3'h6)]))
            begin
              reg295 = reg286;
              reg296 = reg278[(2'h2):(2'h2)];
              reg297 <= (reg279[(2'h2):(1'h0)] ?
                  $signed($unsigned($signed((~reg286)))) : ((reg281 + ("fPglnfCE4gHsa" << reg277)) < wire271));
              reg298 <= ((reg294[(3'h7):(1'h0)] < $unsigned($unsigned(reg294))) >= ((reg279[(2'h3):(1'h0)] ^ {(8'ha5),
                  (wire273 == reg284)}) + ($unsigned(wire272[(2'h2):(1'h1)]) ?
                  reg283[(4'hc):(4'ha)] : reg288[(3'h6):(1'h1)])));
              reg299 = {$unsigned(reg291[(2'h3):(1'h0)])};
            end
          else
            begin
              reg295 <= ($unsigned($signed("H3CZRkBTuP67iwvHf")) < wire271);
              reg296 = $signed($signed((^forvar292[(3'h7):(2'h2)])));
              reg297 = ((reg299[(2'h3):(1'h1)] && (8'ha7)) & ((("MrNmccItsqkLo" > $unsigned((8'had))) ?
                      reg284[(4'h8):(1'h0)] : $unsigned($unsigned((8'h9c)))) ?
                  reg281[(1'h1):(1'h1)] : $unsigned($unsigned(reg281))));
              reg298 <= forvar279[(2'h2):(1'h1)];
            end
          for (forvar300 = (1'h0); (forvar300 < (2'h2)); forvar300 = (forvar300 + (1'h1)))
            begin
              reg301 = (-(!$unsigned((~^wire273[(4'hb):(3'h7)]))));
              reg302 = (!reg288);
              reg303 <= ($signed({(~^$unsigned(reg302)),
                  $unsigned((~wire274))}) >> (8'hbf));
            end
        end
      for (forvar304 = (1'h0); (forvar304 < (2'h2)); forvar304 = (forvar304 + (1'h1)))
        begin
          reg305 = $signed({{{reg281, reg302},
                  ($signed(reg286) || $signed((8'hbd)))}});
          for (forvar306 = (1'h0); (forvar306 < (2'h3)); forvar306 = (forvar306 + (1'h1)))
            begin
              reg307 <= (~{forvar277[(1'h1):(1'h1)]});
              reg308 <= ($signed("8Qs9VmUA55K2JE") >>> reg301);
            end
          if (wire274[(3'h5):(2'h2)])
            begin
              reg309 <= reg293;
              reg310 <= reg290[(3'h5):(3'h4)];
              reg311 <= reg283;
              reg312 = {($unsigned((~|reg311)) ?
                      wire276 : {(wire272[(3'h7):(2'h2)] == (reg278 ?
                              (8'hbe) : reg299)),
                          {{forvar287, reg283}}}),
                  $unsigned($unsigned($signed(reg293)))};
              reg313 <= ((|({reg309} >>> ({reg308} ?
                  ((8'hb2) == (8'hb4)) : $unsigned((8'hbc))))) <<< {reg289[(1'h1):(1'h0)]});
            end
          else
            begin
              reg309 <= ("5S7" * "Vzqn51FqbVrJuW");
              reg310 <= ({reg297[(1'h0):(1'h0)]} - {$unsigned(reg287[(4'hb):(1'h0)]),
                  reg303[(4'hf):(2'h2)]});
              reg311 <= reg277[(3'h5):(2'h2)];
            end
          if (forvar287)
            begin
              reg314 = $unsigned({$unsigned(wire276)});
              reg315 <= forvar287[(3'h4):(2'h3)];
              reg316 <= $signed($unsigned($unsigned(({reg279,
                  reg277} <= ((8'hb0) >>> (8'hac))))));
            end
          else
            begin
              reg314 <= ((|"u5ppwKfFkbF0m") ?
                  (((((8'had) ~^ reg280) ?
                              (forvar300 ^~ reg279) : ((7'h41) <<< reg311)) ?
                          "550xDEyZ0O5MXUElP" : {(8'ha3)}) ?
                      $unsigned(({(8'ha0), forvar304} & (reg315 ?
                          forvar306 : reg302))) : wire274[(1'h0):(1'h0)]) : reg280[(2'h3):(1'h0)]);
              reg315 <= ((reg310 >= forvar277[(1'h1):(1'h1)]) + reg299[(3'h4):(2'h3)]);
              reg316 <= $unsigned((reg283 > $unsigned({(reg296 > (8'hbe))})));
            end
          reg317 <= $signed((reg310 && (wire272 * ($unsigned(reg314) | $signed((8'h9c))))));
        end
      for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
        begin
          for (forvar319 = (1'h0); (forvar319 < (1'h1)); forvar319 = (forvar319 + (1'h1)))
            begin
              reg320 = ((reg317[(3'h6):(3'h6)] ?
                  (^~reg286) : $signed(((wire274 ?
                      reg291 : (8'ha8)) * reg294))) || wire272[(4'h9):(4'h8)]);
            end
          reg321 <= ($signed(wire272[(4'h9):(1'h1)]) < (forvar300 >>> (^(~|$signed(forvar287)))));
          for (forvar322 = (1'h0); (forvar322 < (1'h0)); forvar322 = (forvar322 + (1'h1)))
            begin
              reg323 <= ((8'ha8) > $unsigned(reg296[(2'h3):(2'h3)]));
              reg324 <= (forvar288[(1'h1):(1'h1)] ?
                  (reg277 >> (reg294[(2'h3):(1'h0)] <<< forvar285[(3'h7):(3'h6)])) : wire271[(3'h4):(1'h0)]);
              reg325 <= (reg279 ?
                  ($unsigned($signed((forvar322 > (8'h9f)))) ?
                      $signed(reg302) : {reg307[(5'h13):(4'ha)],
                          (^reg321[(2'h2):(2'h2)])}) : (^({(8'hb8),
                      $unsigned(reg296)} <= ($unsigned((8'ha2)) ?
                      $unsigned((8'ha7)) : reg323))));
            end
          if ($signed((8'hb1)))
            begin
              reg326 = ($unsigned(((reg308 >= {wire274,
                  forvar318}) >> ((reg293 ?
                  reg299 : reg280) - forvar285[(1'h1):(1'h0)]))) ~^ (8'h9f));
              reg327 = (7'h40);
              reg328 <= "mMGOo2GzFOknBGc";
              reg329 <= (7'h42);
            end
          else
            begin
              reg326 = $signed({reg311});
              reg327 <= reg315[(4'ha):(3'h5)];
              reg328 <= ($unsigned((reg290[(4'hc):(3'h7)] ?
                      reg320[(2'h2):(2'h2)] : (8'ha2))) ?
                  (+reg279) : "O5tqTGwS0iRKX4Hn8T");
              reg329 = ("tBsZ4kAtvH1SrCp" ^~ ($unsigned($unsigned({(8'ha4),
                  reg328})) | ((reg280 ?
                  ((8'hae) < (8'had)) : {reg325}) || "UNts0JIXk8sw9")));
              reg330 <= ({{reg321[(3'h5):(2'h2)], wire273}} ?
                  $signed(wire273[(5'h10):(3'h4)]) : (reg308 ?
                      (reg311 ?
                          {reg307} : reg314[(3'h6):(1'h0)]) : $signed({(reg310 ?
                              (8'hb8) : reg312)})));
            end
          for (forvar331 = (1'h0); (forvar331 < (2'h2)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 <= (reg308[(4'ha):(2'h2)] << (($signed($unsigned(forvar287)) > {(|(8'haf)),
                  (reg302 != reg320)}) ^~ ((forvar322[(3'h6):(3'h6)] <= forvar304) <= $signed($signed(forvar285)))));
              reg333 <= ((~^($unsigned($unsigned(reg320)) ?
                  ($signed((8'hb6)) <= ((8'ha6) ?
                      (8'ha0) : reg329)) : {$unsigned(forvar279)})) & (^~forvar304[(4'h9):(3'h6)]));
              reg334 <= $unsigned(($unsigned($signed(reg284)) ?
                  reg283[(3'h6):(3'h4)] : (reg311 < ((|(7'h41)) ^ {reg317,
                      reg284}))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
        begin
          if ((reg326 ?
              reg320[(3'h6):(1'h1)] : (&($unsigned("dv54Ne3BNqh2") + ($unsigned(reg325) || reg277[(4'ha):(2'h2)])))))
            begin
              reg336 = $signed($unsigned(reg320));
              reg337 = ((~^{((^reg316) | {reg290, (8'ha2)}),
                      $unsigned(reg298)}) ?
                  $signed(((~^(reg315 ?
                      forvar285 : reg288)) - (reg301 || (reg324 - forvar292)))) : ($unsigned(wire275) ?
                      ((^(8'ha6)) <= (8'hae)) : reg320));
              reg338 <= $unsigned(($unsigned((7'h40)) && ($unsigned(((8'hae) | reg296)) ?
                  (8'hb2) : (-{reg324, reg329}))));
            end
          else
            begin
              reg336 <= ({"S5yvlf2BYJ"} || reg321);
              reg337 <= ({forvar306[(1'h0):(1'h0)],
                  {$unsigned($unsigned(reg291)),
                      $unsigned(reg303)}} | $unsigned($signed(forvar279)));
              reg338 = $unsigned({$unsigned($unsigned($unsigned((8'hb9))))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg339 = $signed(((^(((7'h43) == reg325) ?
          wire274 : ((7'h43) + forvar306))) + reg329));
      for (forvar340 = (1'h0); (forvar340 < (3'h4)); forvar340 = (forvar340 + (1'h1)))
        begin
          reg341 = (reg299 ~^ $unsigned($unsigned(reg301)));
          for (forvar342 = (1'h0); (forvar342 < (1'h1)); forvar342 = (forvar342 + (1'h1)))
            begin
              reg343 = (((reg302 ?
                  ($signed(wire272) <<< $unsigned(reg324)) : {(8'hb3),
                      reg313}) >= $unsigned(($signed(reg301) ?
                  $unsigned((8'ha0)) : reg312))) | (^~$signed(({reg305,
                  forvar279} != (forvar285 ? reg333 : reg341)))));
              reg344 <= reg329[(1'h0):(1'h0)];
              reg345 <= (7'h44);
              reg346 <= {{$unsigned({reg283})}};
              reg347 <= reg343;
            end
        end
      reg348 = (8'haf);
      reg349 = $signed(reg334[(2'h3):(1'h1)]);
      reg350 <= (forvar342 ~^ (^$signed((reg288[(4'he):(1'h1)] >>> {reg343}))));
    end
  always
    @(posedge clk) begin
      if ({{$signed(($unsigned(reg334) ^ (7'h40)))},
          $unsigned(($signed($unsigned(forvar277)) <= $unsigned((forvar306 >>> (7'h43)))))})
        begin
          reg351 = $unsigned({{(reg284 << ((7'h40) ^ reg346)), forvar331}});
          for (forvar352 = (1'h0); (forvar352 < (2'h2)); forvar352 = (forvar352 + (1'h1)))
            begin
              reg353 <= {reg283[(4'hc):(4'hb)], "Sruf6tX99cRwSZLdzS4"};
              reg354 <= reg303;
            end
          reg355 <= (({((reg310 ? reg343 : (8'hbe)) ~^ (7'h42)),
              (reg291[(4'h8):(1'h0)] ?
                  ((7'h41) ? (8'hbb) : reg345) : (reg278 ?
                      (8'hb5) : wire273))} >>> reg350) ^~ $unsigned(reg303));
          reg356 <= ($unsigned(($signed({reg310}) != ((wire272 ?
                  reg311 : forvar300) ?
              $signed(reg282) : {reg315}))) - (~^"Pt5UAGnnLBwYfl6ViJN4"));
        end
      else
        begin
          for (forvar351 = (1'h0); (forvar351 < (1'h1)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 <= $unsigned((^reg316));
              reg353 = ((reg288 || reg294) * reg330);
              reg354 <= (|(~wire273));
              reg355 = ({$unsigned($signed($unsigned(reg311)))} && $signed({(reg330[(4'hd):(2'h3)] ^~ forvar318)}));
              reg356 <= $signed(((reg332 == (reg298[(4'h8):(2'h3)] ?
                      reg328 : wire273[(4'hd):(3'h6)])) ?
                  (reg313[(3'h4):(2'h2)] | {forvar304[(3'h6):(1'h0)],
                      $unsigned(forvar335)}) : reg326[(3'h6):(3'h5)]));
            end
          for (forvar357 = (1'h0); (forvar357 < (3'h4)); forvar357 = (forvar357 + (1'h1)))
            begin
              reg358 <= reg307[(5'h12):(4'hb)];
              reg359 <= (reg338[(2'h2):(2'h2)] ?
                  (|{reg312}) : {$unsigned((reg321 ?
                          (reg288 || (8'h9d)) : (~|(8'ha2))))});
            end
          reg360 = {$unsigned({$signed({reg350})})};
          reg361 <= ($unsigned(("3qvQvWBss66xotdw" * reg332[(3'h5):(3'h4)])) && {({$unsigned(reg315)} ?
                  $unsigned((8'ha2)) : $unsigned($signed((8'hb2))))});
        end
    end
  always
    @(posedge clk) begin
      reg362 <= reg311;
      reg363 = (^~$unsigned((8'hab)));
      reg364 <= reg298[(3'h7):(3'h6)];
      for (forvar365 = (1'h0); (forvar365 < (2'h2)); forvar365 = (forvar365 + (1'h1)))
        begin
          for (forvar366 = (1'h0); (forvar366 < (2'h2)); forvar366 = (forvar366 + (1'h1)))
            begin
              reg367 <= (7'h42);
            end
          reg368 = {$unsigned(({reg296,
                  ((8'ha4) <= (8'hbf))} <<< $signed(((7'h41) << reg328)))),
              $unsigned(reg298[(4'ha):(3'h4)])};
        end
      reg369 <= ($signed({$unsigned($unsigned(reg347)),
          $unsigned(((7'h44) >= wire274))}) && ($signed(reg363[(3'h6):(3'h4)]) | forvar342[(2'h3):(1'h1)]));
    end
  always
    @(posedge clk) begin
      if (({({$signed(forvar292), {(8'ha8), (8'hbe)}} ?
              (~&$unsigned(reg344)) : $signed(reg280[(1'h0):(1'h0)])),
          (forvar306[(4'h9):(2'h3)] ?
              reg307 : (8'hbe))} >= ("d1krpw" >>> ({$unsigned(reg333),
              $unsigned(reg346)} ?
          $signed({(8'had), (8'ha2)}) : ((wire273 ? reg297 : reg332) ?
              $unsigned((8'ha5)) : (reg298 ? reg284 : forvar288))))))
        begin
          for (forvar370 = (1'h0); (forvar370 < (1'h1)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 <= ((("f" ?
                  "Yf8ve3" : reg362) || $unsigned($signed({reg346,
                  reg344}))) && ((+($unsigned(reg309) ? reg294 : (~^reg283))) ?
                  $unsigned(reg360) : (reg316[(3'h4):(2'h3)] - {(&reg316),
                      reg352})));
            end
          for (forvar372 = (1'h0); (forvar372 < (1'h1)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 <= ((8'hb9) + {reg303[(3'h4):(2'h3)], reg284});
              reg374 <= $signed((8'hbf));
              reg375 <= ((-reg316[(2'h3):(1'h0)]) ^ reg288);
            end
          reg376 = {reg361[(4'h8):(1'h0)],
              ({$unsigned($unsigned((8'hba)))} ?
                  reg352[(1'h1):(1'h0)] : $unsigned($unsigned($unsigned(reg344))))};
          for (forvar377 = (1'h0); (forvar377 < (3'h4)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 <= {((((reg314 ~^ forvar277) ?
                          $signed((8'hb7)) : $signed((7'h42))) ?
                      ((reg363 <<< reg321) < (reg355 >>> reg315)) : $signed((-reg313))) >= (~&reg329[(2'h2):(1'h1)]))};
              reg379 <= {reg309[(3'h4):(2'h2)]};
              reg380 = {(&((8'haa) ?
                      $unsigned(reg316) : reg368[(4'hc):(4'hc)])),
                  {(+$signed((reg356 + forvar365)))}};
              reg381 <= $unsigned($signed(forvar365[(1'h1):(1'h0)]));
            end
          reg382 <= {$signed(($unsigned("") >> ((reg349 ^ (8'hac)) ?
                  ((8'hbb) || (8'hbd)) : ((8'hb3) >> (8'h9d))))),
              reg349[(1'h1):(1'h1)]};
        end
      else
        begin
          if (reg282)
            begin
              reg370 <= reg362[(4'hf):(4'hd)];
            end
          else
            begin
              reg370 <= reg312[(3'h7):(2'h3)];
              reg371 <= (&reg350[(3'h4):(1'h1)]);
              reg372 <= $unsigned($unsigned(((!"Dp6vJtU7J7EIgdkT6c") >>> forvar288[(4'hb):(1'h0)])));
              reg373 = ($unsigned({$unsigned({forvar340, reg333}),
                  forvar285[(1'h0):(1'h0)]}) == $signed(reg347));
              reg374 = reg311;
            end
          reg375 <= (^~((8'hb1) ?
              $unsigned((reg291 ?
                  (reg341 < reg339) : {reg279,
                      wire271})) : reg277[(4'ha):(3'h4)]));
          reg376 = (reg361 ^~ $signed($unsigned((8'hab))));
        end
      reg383 <= reg296;
    end
  assign wire384 = {reg337[(2'h3):(1'h1)]};
  assign wire385 = $unsigned(reg370);
  assign wire386 = (reg315 >>> reg329[(4'h8):(3'h6)]);
  always
    @(posedge clk) begin
      if ({(8'ha7)})
        begin
          if (reg363)
            begin
              reg387 <= (reg311 & wire271[(4'ha):(2'h3)]);
              reg388 = (~$unsigned($unsigned(reg338[(2'h2):(1'h1)])));
              reg389 <= (7'h43);
              reg390 = ({"1PeRENi", forvar285} == ({$unsigned({reg375,
                      (7'h40)})} ^~ (~|reg302[(3'h6):(3'h6)])));
              reg391 <= $unsigned({$unsigned(reg380),
                  forvar300[(1'h0):(1'h0)]});
            end
          else
            begin
              reg387 = (reg351 >>> (^~reg380));
              reg388 = (reg308 && (&((&{reg303}) ?
                  $unsigned({(8'hae)}) : (((8'hb7) >= reg371) == (~forvar300)))));
              reg389 <= reg360[(3'h4):(2'h2)];
              reg390 <= (reg315 ?
                  (-{{(~|reg389)}}) : {wire271[(3'h7):(3'h5)], "SPJx"});
            end
          reg392 <= $unsigned("MJEyCxNOGYV");
          for (forvar393 = (1'h0); (forvar393 < (1'h0)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= ((8'hbb) + (reg281 ?
                  ((reg310[(1'h0):(1'h0)] != (forvar306 >= wire274)) == ({(8'hbe),
                          reg334} ?
                      reg284[(4'hb):(4'h8)] : forvar352)) : $unsigned(reg293)));
              reg395 = "bTXQdoHR";
              reg396 <= $signed(reg280);
            end
          if ((|(reg383[(1'h1):(1'h0)] << reg396)))
            begin
              reg397 <= (+(reg328 != $unsigned((+reg372[(3'h4):(1'h1)]))));
              reg398 = ($unsigned({$unsigned(((8'ha8) ? reg290 : wire271))}) ?
                  ((($unsigned((8'ha3)) ?
                          (7'h40) : ((8'ha7) >>> reg332)) >>> ($unsigned(reg293) ^ {forvar318})) ?
                      wire272 : (~^{reg394})) : {reg314[(2'h3):(1'h1)],
                      {(forvar351[(4'h9):(3'h4)] < ((8'ha0) * reg352))}});
            end
          else
            begin
              reg397 = $unsigned(($unsigned($unsigned((8'hbb))) <<< $signed(reg363[(3'h4):(2'h2)])));
              reg398 <= $unsigned(reg336[(4'hb):(3'h6)]);
              reg399 <= reg388[(4'hf):(4'ha)];
              reg400 <= forvar285[(1'h1):(1'h0)];
              reg401 <= "UeGxkClYHm6RKN0";
            end
          reg402 <= $unsigned($unsigned({(8'hbe),
              $unsigned({reg320, reg369})}));
        end
      else
        begin
          reg387 = (~($signed(((reg287 > reg345) ?
              $signed(forvar342) : reg397[(4'he):(2'h3)])) == reg370[(2'h3):(1'h1)]));
          for (forvar388 = (1'h0); (forvar388 < (2'h3)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 <= {$signed({((reg383 && reg368) != "O0p4U1xlKoV"),
                      (8'hab)})};
              reg390 <= $unsigned($signed(reg282));
              reg391 <= ($unsigned({$unsigned({(8'haf), reg389}),
                  ((reg337 && forvar366) + $unsigned(reg390))}) && {$unsigned({reg339[(3'h4):(1'h0)]}),
                  (reg294[(1'h0):(1'h0)] + $unsigned((forvar322 ?
                      reg396 : forvar304)))});
              reg392 <= $unsigned((8'ha8));
            end
          for (forvar393 = (1'h0); (forvar393 < (1'h0)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 = (~&reg298);
              reg395 <= (reg279 != (8'had));
            end
          reg396 <= $signed((~&forvar287[(3'h4):(2'h2)]));
          reg397 = ({(((&(8'hbb)) ? reg315[(4'ha):(3'h5)] : (~reg321)) ?
                  forvar318 : $unsigned((reg352 || (8'hb9))))} >> reg387[(2'h2):(1'h1)]);
        end
      if ("k3wRrh6XNiky9FulHI")
        begin
          for (forvar403 = (1'h0); (forvar403 < (1'h1)); forvar403 = (forvar403 + (1'h1)))
            begin
              reg404 = $unsigned($unsigned({{((8'hbf) ? reg400 : reg395)}}));
            end
          reg405 = {wire386};
          reg406 <= (~|(&(8'ha7)));
          for (forvar407 = (1'h0); (forvar407 < (1'h0)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 <= $signed({$unsigned(((reg308 ?
                      (8'ha1) : (8'hae)) ^~ forvar366[(2'h2):(1'h1)])),
                  (reg294 <= {reg338[(1'h0):(1'h0)],
                      (reg310 ? reg337 : reg347)})});
              reg409 = ((|reg309) && ({reg351,
                  $unsigned(reg280)} >>> reg341[(4'hc):(3'h5)]));
              reg410 <= $signed((forvar322[(3'h7):(2'h3)] ?
                  (&$unsigned(reg395[(3'h4):(2'h2)])) : reg405));
              reg411 = $unsigned((reg311 - $unsigned($signed((8'h9f)))));
            end
          reg412 <= reg400[(2'h2):(1'h1)];
        end
      else
        begin
          reg403 <= ($signed("5txM1rA4") + $unsigned(reg307));
          reg404 = ((&{forvar318}) ~^ $signed($unsigned((8'hb1))));
          for (forvar405 = (1'h0); (forvar405 < (2'h3)); forvar405 = (forvar405 + (1'h1)))
            begin
              reg406 <= {$unsigned((~^($unsigned(reg333) ?
                      (!wire385) : (reg308 && forvar342)))),
                  (+$unsigned(forvar340[(2'h3):(2'h3)]))};
              reg407 = $unsigned({"MD8d4qpqU",
                  (forvar292 >> $signed($signed(forvar357)))});
            end
        end
      reg413 = reg332[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg414 <= ($signed($signed(reg358[(4'hc):(3'h6)])) || $unsigned($unsigned(((!forvar352) > forvar351[(3'h4):(2'h2)]))));
      reg415 <= forvar351[(3'h7):(1'h1)];
      reg416 = (&forvar335[(2'h2):(2'h2)]);
      reg417 <= $unsigned(($signed($signed($signed(reg396))) ?
          reg330 : {{$unsigned(reg363)}}));
      for (forvar418 = (1'h0); (forvar418 < (1'h1)); forvar418 = (forvar418 + (1'h1)))
        begin
          for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 <= {wire272, reg349};
              reg421 <= reg288[(4'hb):(4'h8)];
              reg422 = (forvar407[(1'h0):(1'h0)] ?
                  reg382[(3'h4):(3'h4)] : $unsigned(reg403[(2'h2):(1'h1)]));
              reg423 <= ((-{reg391[(4'h8):(1'h1)],
                  {wire385[(3'h5):(1'h0)]}}) <<< $unsigned(($unsigned((forvar357 ^~ (8'ha8))) >>> $unsigned(reg402[(1'h0):(1'h0)]))));
              reg424 <= $signed(((8'hb2) ?
                  {(reg410 != {(8'ha2)}),
                      {reg328[(4'hb):(1'h1)]}} : $unsigned(($unsigned(reg346) >= reg287[(4'h9):(3'h6)]))));
            end
          for (forvar425 = (1'h0); (forvar425 < (3'h4)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 = (^reg284[(4'he):(3'h7)]);
              reg427 = ($unsigned(((reg396[(1'h0):(1'h0)] <= reg313[(3'h7):(1'h0)]) ?
                      reg353 : $signed(((8'hb1) ? reg281 : reg355)))) ?
                  reg359[(1'h0):(1'h0)] : $unsigned($signed(($unsigned(forvar300) | $unsigned(forvar388)))));
              reg428 <= $unsigned(reg427[(4'h8):(3'h7)]);
              reg429 <= (($unsigned(reg376[(2'h2):(2'h2)]) ?
                      forvar319[(1'h1):(1'h1)] : ((reg323 != reg325) + (reg305 + reg328))) ?
                  {reg345,
                      (reg327 != (~|$signed((8'ha3))))} : ({(forvar300 >= (&reg390)),
                          $unsigned((forvar304 >>> forvar285))} ?
                      (reg378 ? reg410 : reg297) : {$signed(reg374)}));
              reg430 <= reg280;
            end
          for (forvar431 = (1'h0); (forvar431 < (2'h3)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 <= $signed(("2u5B9UnFyM" ?
                  (8'ha8) : ((&$unsigned((8'hab))) ?
                      $signed($unsigned((7'h41))) : ($unsigned(reg294) << reg405[(1'h0):(1'h0)]))));
              reg433 = (($unsigned(((reg324 * forvar405) ?
                      (forvar365 ?
                          reg279 : reg348) : (forvar393 * reg427))) != reg347[(2'h2):(1'h0)]) ?
                  (|{(8'had),
                      (8'hb9)}) : $unsigned($signed($unsigned({reg409}))));
              reg434 <= {(^(~&reg287)), reg368};
            end
          reg435 = {(8'h9c)};
          if ($unsigned(reg320))
            begin
              reg436 <= $signed($unsigned($unsigned(wire272)));
              reg437 <= ((((7'h40) - $signed({reg311,
                  reg435})) == reg396) != $signed((reg297 < $unsigned(reg436[(4'ha):(3'h5)]))));
              reg438 <= (((!{{reg289},
                  reg378[(3'h7):(3'h7)]}) == (-forvar331[(3'h5):(1'h1)])) && $signed((-(|$unsigned(reg324)))));
              reg439 = $signed(reg391[(2'h2):(2'h2)]);
              reg440 = reg370[(4'hb):(3'h7)];
            end
          else
            begin
              reg436 <= ((($signed((8'hb7)) ?
                          (^~$unsigned(reg401)) : (-(forvar357 ?
                              (8'h9e) : reg333))) ?
                      reg415 : (~^(reg290[(4'hd):(4'ha)] > reg278))) ?
                  (($signed(reg361) ?
                      reg329[(3'h5):(1'h1)] : (forvar319 ^ "2MO8VTgP")) ^ ($unsigned($signed(reg396)) && ($unsigned((8'hb0)) ?
                      $unsigned(reg297) : (reg294 ?
                          reg436 : reg367)))) : (reg334 != ((~$unsigned(forvar342)) < reg281[(1'h1):(1'h0)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg441 <= (({(&(~|(8'ha0))), $signed(forvar322)} & reg395) ?
          $unsigned(reg403[(4'h8):(2'h2)]) : reg412[(1'h1):(1'h0)]);
      reg442 = ((8'hae) << $unsigned({($signed(reg376) + $signed(reg417)),
          ((8'hbe) && (8'hb0))}));
    end
  always
    @(posedge clk) begin
      if (reg294[(1'h0):(1'h0)])
        begin
          reg443 <= $unsigned((((^$unsigned((8'ha0))) ? {forvar331} : "qyJWl") ?
              {{(~forvar285),
                      $unsigned(reg364)}} : $unsigned(((reg317 ~^ reg404) ?
                  {(8'ha2)} : (8'ha6)))));
          for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 = $signed($unsigned((8'hb1)));
              reg446 <= (8'h9c);
              reg447 = $unsigned(wire271[(3'h4):(1'h0)]);
              reg448 = (&((8'h9c) < reg344[(1'h1):(1'h0)]));
            end
        end
      else
        begin
          reg443 <= wire271[(4'hb):(1'h0)];
          reg444 <= reg287[(3'h4):(1'h0)];
          reg445 <= {$unsigned((+((reg421 ? (8'ha6) : reg326) ^~ ((8'ha5) ?
                  (7'h43) : reg387)))),
              (reg311 >= $signed(reg354))};
          reg446 = "DrN8";
        end
      reg449 <= reg356;
    end
  assign wire450 = {"Z"};
  assign wire451 = reg301;
  always
    @(posedge clk) begin
      for (forvar452 = (1'h0); (forvar452 < (3'h4)); forvar452 = (forvar452 + (1'h1)))
        begin
          reg453 <= reg363;
          reg454 = {reg442[(4'hd):(3'h6)],
              {($unsigned($unsigned((8'hbd))) & (reg321[(4'hc):(4'h9)] * reg367[(3'h4):(2'h2)]))}};
          for (forvar455 = (1'h0); (forvar455 < (2'h2)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 <= wire385;
              reg457 <= reg401[(2'h3):(1'h1)];
            end
          reg458 <= reg290;
          for (forvar459 = (1'h0); (forvar459 < (2'h3)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 = reg277;
              reg461 <= forvar340;
              reg462 <= (forvar455[(2'h3):(1'h0)] >>> $signed(forvar459[(3'h5):(1'h1)]));
              reg463 <= $unsigned($signed(reg408[(1'h1):(1'h1)]));
              reg464 = {(reg421[(3'h7):(3'h5)] ?
                      ((8'hae) ?
                          forvar370 : ({reg416,
                              (8'ha5)} & (8'hbf))) : (!reg341)),
                  ({(reg429 ?
                          (8'ha8) : (reg407 ?
                              (8'hb9) : (8'h9f)))} || reg440[(3'h4):(2'h2)])};
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar465 = (1'h0); (forvar465 < (1'h1)); forvar465 = (forvar465 + (1'h1)))
        begin
          if ((($signed((+(forvar300 ~^ reg426))) < (reg324 ^ (!$signed(reg427)))) == $unsigned(((((8'hbe) ?
              reg286 : forvar419) && $signed(reg281)) - (8'ha3)))))
            begin
              reg466 <= $unsigned(({(reg413 ?
                          reg321[(4'h9):(4'h8)] : $unsigned(reg354))} ?
                  (reg303[(5'h10):(2'h3)] ?
                      (8'hb9) : $unsigned((~^reg317))) : (8'ha2)));
              reg467 <= forvar331[(3'h5):(3'h5)];
              reg468 <= (((!$unsigned((reg414 | reg372))) ?
                  forvar365 : $unsigned($unsigned({(8'ha4)}))) > forvar403[(3'h5):(3'h5)]);
              reg469 <= forvar370[(4'h9):(3'h6)];
            end
          else
            begin
              reg466 <= {{{(reg414 ? "X3Ysfz" : reg280)}},
                  ({((reg281 ? reg389 : reg370) ?
                          (8'ha1) : $unsigned(reg411))} && reg449[(4'ha):(3'h6)])};
              reg467 = {$signed((8'hbb)), (~^{reg291[(2'h3):(2'h2)]})};
              reg468 <= (($signed(((8'hbd) <= (reg355 == reg312))) >> ($unsigned(reg277) >> {{wire385}})) >>> reg398);
              reg469 <= {(+(!(8'hb6)))};
            end
          for (forvar470 = (1'h0); (forvar470 < (3'h4)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 = {($unsigned(reg345[(2'h2):(1'h1)]) + $unsigned(reg345))};
              reg472 = (reg326 ~^ reg317);
              reg473 <= reg352[(4'hc):(4'h8)];
            end
        end
      reg474 = {$unsigned($unsigned(wire450[(1'h1):(1'h1)])), (~|reg362)};
    end
  assign wire475 = {$signed(((8'hb8) && wire384[(4'hc):(3'h6)]))};
  always
    @(posedge clk) begin
      if (forvar287[(3'h4):(2'h2)])
        begin
          reg476 = ((reg443 + (~|{(~|forvar393),
              (8'haa)})) - (wire475[(3'h4):(3'h4)] == {((reg368 >= reg372) ?
                  $unsigned(reg412) : reg286[(1'h0):(1'h0)]),
              reg391}));
        end
      else
        begin
          reg476 <= $unsigned(reg443);
          reg477 <= $unsigned(reg416[(3'h4):(3'h4)]);
          reg478 = ($signed($unsigned((reg320[(4'h8):(4'h8)] == $signed((8'hba))))) >= reg416);
          reg479 <= ($unsigned((^~(reg415[(1'h1):(1'h1)] ~^ (wire386 ^~ reg436)))) ?
              ((!$signed(((8'ha0) ?
                  reg310 : reg401))) ^ (reg296[(4'ha):(4'h9)] ?
                  $unsigned((reg283 ? forvar407 : (8'h9e))) : (^((8'ha2) ?
                      reg332 : forvar300)))) : (8'ha5));
          for (forvar480 = (1'h0); (forvar480 < (2'h3)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= ({$signed((reg343 > $unsigned(forvar370))),
                  (((~|(8'hbb)) ? (7'h42) : reg324[(2'h2):(1'h1)]) * ((8'haf) ?
                      reg368 : $signed(reg435)))} & (reg427[(3'h7):(2'h3)] ?
                  ($unsigned($unsigned((8'hb4))) ?
                      $unsigned({reg293,
                          (8'ha2)}) : reg473[(2'h3):(2'h2)]) : reg307));
              reg482 = wire271[(4'h8):(2'h2)];
              reg483 <= (reg328[(3'h6):(3'h4)] & {$unsigned(((forvar331 ?
                          reg460 : reg348) ?
                      (reg390 <<< reg309) : (reg407 ? (8'ha1) : (7'h42)))),
                  (forvar405 <= (reg461[(2'h3):(2'h2)] ^~ {(7'h43), reg332}))});
              reg484 <= (reg430[(2'h3):(1'h0)] + (8'ha3));
              reg485 <= (8'ha2);
            end
        end
      for (forvar486 = (1'h0); (forvar486 < (1'h1)); forvar486 = (forvar486 + (1'h1)))
        begin
          reg487 <= forvar279[(4'h8):(2'h3)];
          if ($unsigned(reg401[(1'h0):(1'h0)]))
            begin
              reg488 <= reg370[(4'hc):(2'h3)];
              reg489 = (^~$unsigned({reg371, reg356}));
              reg490 <= ({(reg310 ? reg473 : (8'hba)),
                      ("VyZg" ?
                          $unsigned($unsigned(reg469)) : $signed((reg395 ?
                              reg422 : forvar306)))} ?
                  reg325 : ({{(forvar372 ? reg286 : (8'haf))},
                      {reg278, (-reg369)}} && $signed({forvar388[(4'hb):(4'h8)],
                      reg362[(4'hc):(4'hc)]})));
            end
          else
            begin
              reg488 = reg397;
              reg489 <= {$unsigned($unsigned($unsigned($signed(forvar285)))),
                  (reg282[(2'h3):(2'h3)] & (&("pImPydzTNOIULo" ?
                      $unsigned((8'hb1)) : {(8'haf)})))};
            end
          reg491 <= ({$signed($signed(reg345))} >>> (forvar470[(3'h6):(3'h5)] == (^(~|reg315[(4'h8):(3'h7)]))));
          reg492 = (~^reg324);
          reg493 <= (($signed($unsigned($unsigned(forvar365))) ?
              reg360[(3'h7):(3'h5)] : forvar352) || (&($unsigned((~reg403)) | ($unsigned(reg481) ^~ $signed(reg438)))));
        end
      reg494 <= (8'hbd);
      for (forvar495 = (1'h0); (forvar495 < (1'h0)); forvar495 = (forvar495 + (1'h1)))
        begin
          if ((reg442[(3'h5):(1'h0)] * (8'ha8)))
            begin
              reg496 <= (8'hb7);
            end
          else
            begin
              reg496 <= (7'h42);
              reg497 <= reg337[(3'h4):(1'h1)];
            end
          for (forvar498 = (1'h0); (forvar498 < (2'h3)); forvar498 = (forvar498 + (1'h1)))
            begin
              reg499 = forvar405;
              reg500 = (reg461[(1'h1):(1'h1)] <<< $unsigned($unsigned(forvar455[(1'h0):(1'h0)])));
              reg501 <= forvar288[(4'ha):(3'h6)];
              reg502 = wire272[(3'h5):(3'h5)];
            end
        end
      for (forvar503 = (1'h0); (forvar503 < (1'h0)); forvar503 = (forvar503 + (1'h1)))
        begin
          reg504 <= ($unsigned(($signed((8'ha6)) - reg435)) * forvar403);
          reg505 <= $unsigned({reg396});
          for (forvar506 = (1'h0); (forvar506 < (1'h1)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 = (($unsigned(((reg445 <<< forvar388) == reg412[(1'h0):(1'h0)])) ?
                  {$unsigned({forvar352}),
                      {$signed(reg349)}} : reg484[(4'h9):(3'h6)]) >>> (($signed($unsigned(forvar366)) * ((reg355 >= (8'hb4)) << {forvar470,
                      (8'hae)})) ?
                  {(8'ha4)} : {forvar342}));
              reg508 = (reg445 ?
                  {"YT0DR51"} : $unsigned((($unsigned(reg440) ^~ {reg293,
                      (8'hb5)}) >> reg295)));
              reg509 <= (8'hb6);
            end
        end
    end
  assign wire510 = ($signed(forvar425) < reg405[(4'hc):(4'hc)]);
  assign wire511 = forvar372[(2'h2):(1'h0)];
  assign wire512 = forvar419;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module109
#( parameter param266 = (^~(!((((8'ha2) | (8'hb3)) - ((8'ha0) >> (8'hbd))) ^ {((8'hac) && (8'hbb))})))
, parameter param267 = param266 )
(y, clk, wire114, wire113, wire112, wire111, wire110);
  output wire [(32'h74e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire114;
  input wire [(4'hb):(1'h0)] wire113;
  input wire [(4'hc):(1'h0)] wire112;
  input wire [(5'h12):(1'h0)] wire111;
  input wire signed [(5'h12):(1'h0)] wire110;
  wire [(4'h8):(1'h0)] wire265;
  wire signed [(5'h15):(1'h0)] wire264;
  wire signed [(5'h13):(1'h0)] wire263;
  wire signed [(5'h15):(1'h0)] wire262;
  wire signed [(4'hd):(1'h0)] wire261;
  wire [(3'h5):(1'h0)] wire260;
  reg [(2'h3):(1'h0)] reg259 = (1'h0);
  reg [(4'h8):(1'h0)] reg258 = (1'h0);
  reg [(3'h7):(1'h0)] reg257 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg256 = (1'h0);
  reg [(3'h4):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar253 = (1'h0);
  reg signed [(4'he):(1'h0)] reg252 = (1'h0);
  reg [(4'he):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg250 = (1'h0);
  reg [(5'h13):(1'h0)] forvar249 = (1'h0);
  reg [(4'hb):(1'h0)] forvar248 = (1'h0);
  reg [(5'h12):(1'h0)] reg247 = (1'h0);
  reg [(3'h6):(1'h0)] forvar246 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg245 = (1'h0);
  reg [(4'he):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar243 = (1'h0);
  reg [(5'h12):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg241 = (1'h0);
  reg [(3'h6):(1'h0)] forvar239 = (1'h0);
  reg [(4'hf):(1'h0)] forvar236 = (1'h0);
  reg [(4'h9):(1'h0)] reg234 = (1'h0);
  reg [(5'h11):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg236 = (1'h0);
  reg [(5'h11):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar234 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg233 = (1'h0);
  reg [(2'h3):(1'h0)] reg232 = (1'h0);
  wire [(4'he):(1'h0)] wire231;
  wire [(4'hb):(1'h0)] wire230;
  wire signed [(5'h12):(1'h0)] wire229;
  wire signed [(2'h3):(1'h0)] wire228;
  reg signed [(3'h5):(1'h0)] reg227 = (1'h0);
  reg [(5'h14):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg225 = (1'h0);
  reg [(4'h8):(1'h0)] reg224 = (1'h0);
  reg [(2'h2):(1'h0)] reg223 = (1'h0);
  reg [(4'h8):(1'h0)] reg222 = (1'h0);
  reg [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg220 = (1'h0);
  reg [(3'h5):(1'h0)] forvar219 = (1'h0);
  reg [(3'h6):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg217 = (1'h0);
  reg [(5'h13):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg215 = (1'h0);
  reg [(4'hf):(1'h0)] reg214 = (1'h0);
  reg [(2'h2):(1'h0)] reg213 = (1'h0);
  wire [(4'hb):(1'h0)] wire212;
  reg signed [(4'h9):(1'h0)] reg211 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar210 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg209 = (1'h0);
  reg [(2'h3):(1'h0)] reg208 = (1'h0);
  reg [(5'h14):(1'h0)] reg207 = (1'h0);
  reg [(5'h12):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar205 = (1'h0);
  reg [(4'h8):(1'h0)] reg204 = (1'h0);
  reg [(5'h14):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg [(5'h13):(1'h0)] reg201 = (1'h0);
  reg [(5'h11):(1'h0)] forvar200 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg198 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg197 = (1'h0);
  reg [(4'hf):(1'h0)] reg196 = (1'h0);
  reg [(5'h12):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg194 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar193 = (1'h0);
  reg [(2'h3):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg191 = (1'h0);
  reg [(4'hb):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg189 = (1'h0);
  reg [(2'h3):(1'h0)] reg188 = (1'h0);
  reg [(4'hb):(1'h0)] reg187 = (1'h0);
  reg [(5'h13):(1'h0)] reg186 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar185 = (1'h0);
  reg [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(2'h2):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg182 = (1'h0);
  reg [(5'h15):(1'h0)] reg181 = (1'h0);
  reg [(4'hc):(1'h0)] forvar180 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg179 = (1'h0);
  reg [(4'h9):(1'h0)] reg178 = (1'h0);
  reg [(4'hc):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg176 = (1'h0);
  reg [(2'h2):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg174 = (1'h0);
  reg signed [(4'he):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg170 = (1'h0);
  reg [(5'h14):(1'h0)] reg169 = (1'h0);
  reg [(4'h8):(1'h0)] forvar168 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg164 = (1'h0);
  reg [(2'h2):(1'h0)] reg163 = (1'h0);
  reg [(4'hd):(1'h0)] reg162 = (1'h0);
  reg [(4'ha):(1'h0)] reg161 = (1'h0);
  reg [(5'h15):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] forvar153 = (1'h0);
  reg [(3'h7):(1'h0)] reg152 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg156 = (1'h0);
  reg [(5'h15):(1'h0)] reg155 = (1'h0);
  reg [(3'h5):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg153 = (1'h0);
  reg [(3'h6):(1'h0)] forvar152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar149 = (1'h0);
  reg [(3'h4):(1'h0)] reg139 = (1'h0);
  reg [(5'h11):(1'h0)] reg148 = (1'h0);
  reg [(3'h4):(1'h0)] reg147 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg144 = (1'h0);
  reg [(3'h6):(1'h0)] forvar143 = (1'h0);
  reg [(4'hc):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg141 = (1'h0);
  reg [(4'ha):(1'h0)] reg140 = (1'h0);
  reg [(5'h14):(1'h0)] forvar139 = (1'h0);
  reg [(4'hf):(1'h0)] reg138 = (1'h0);
  wire [(4'hb):(1'h0)] wire137;
  wire [(4'hf):(1'h0)] wire136;
  wire [(4'h9):(1'h0)] wire135;
  reg [(3'h4):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg132 = (1'h0);
  reg [(4'he):(1'h0)] reg131 = (1'h0);
  reg [(4'hf):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg129 = (1'h0);
  reg [(3'h4):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg127 = (1'h0);
  reg [(2'h3):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar125 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] reg122 = (1'h0);
  reg [(2'h2):(1'h0)] reg121 = (1'h0);
  reg [(5'h11):(1'h0)] reg120 = (1'h0);
  reg [(3'h5):(1'h0)] forvar119 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg [(4'hf):(1'h0)] forvar116 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg115 = (1'h0);
  assign y = {wire265,
                 wire264,
                 wire263,
                 wire262,
                 wire261,
                 wire260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 forvar253,
                 reg252,
                 reg251,
                 reg250,
                 forvar249,
                 forvar248,
                 reg247,
                 forvar246,
                 reg245,
                 reg244,
                 forvar243,
                 reg242,
                 reg241,
                 forvar239,
                 forvar236,
                 reg234,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 forvar234,
                 reg233,
                 reg232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 wire212,
                 reg211,
                 forvar210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 forvar205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 forvar200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 forvar193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 forvar185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 forvar180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 forvar168,
                 forvar164,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 forvar158,
                 reg157,
                 forvar153,
                 reg152,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 forvar152,
                 reg151,
                 reg150,
                 forvar149,
                 reg139,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 reg141,
                 reg140,
                 forvar139,
                 reg138,
                 wire137,
                 wire136,
                 wire135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 forvar125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 forvar119,
                 reg118,
                 reg117,
                 forvar116,
                 reg115,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg115 <= $unsigned((~|({$signed(wire112),
          (wire112 << wire110)} < ((wire113 >= (8'ha3)) <= $signed((8'hbe))))));
      for (forvar116 = (1'h0); (forvar116 < (2'h2)); forvar116 = (forvar116 + (1'h1)))
        begin
          reg117 <= {wire110};
          reg118 = {reg115};
          for (forvar119 = (1'h0); (forvar119 < (3'h4)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 <= ({wire113[(3'h7):(3'h5)]} != reg118);
              reg121 <= (~((($unsigned(reg115) ?
                      (reg118 ? reg115 : (7'h41)) : {(8'h9c), wire112}) ?
                  forvar119[(1'h0):(1'h0)] : {reg117[(4'h9):(1'h1)],
                      wire114[(1'h1):(1'h0)]}) & ((~&(^(8'h9d))) ?
                  $unsigned((^(8'hac))) : wire110[(4'h9):(3'h4)])));
              reg122 = wire112[(2'h2):(1'h0)];
              reg123 = ($unsigned(wire113[(4'h8):(3'h6)]) ?
                  reg117 : $signed(reg117[(3'h4):(1'h1)]));
              reg124 <= (8'h9f);
            end
          for (forvar125 = (1'h0); (forvar125 < (2'h3)); forvar125 = (forvar125 + (1'h1)))
            begin
              reg126 <= forvar119;
              reg127 <= $signed($signed($unsigned((wire111[(5'h10):(3'h6)] ?
                  $unsigned(reg115) : {(8'ha2), wire114}))));
              reg128 <= ((~&(8'ha2)) || wire114[(2'h2):(1'h1)]);
              reg129 <= reg128;
              reg130 = $unsigned(reg121[(2'h2):(1'h1)]);
            end
          if ((forvar116 ?
              $signed(reg120[(5'h10):(3'h6)]) : (!(wire110 <<< ((~&(8'hbc)) ?
                  (reg129 ? reg122 : reg117) : forvar116[(4'ha):(3'h6)])))))
            begin
              reg131 = reg120;
              reg132 = reg121[(1'h1):(1'h0)];
              reg133 = ($signed((((forvar125 == (8'ha3)) != $unsigned(reg131)) ?
                  ({reg122} ^~ reg118) : ({forvar125} == reg132))) != reg120[(2'h2):(1'h0)]);
            end
          else
            begin
              reg131 = {(($unsigned((reg120 == (8'ha0))) ?
                      $unsigned((forvar116 | (8'ha8))) : reg121[(2'h2):(1'h1)]) + reg121[(1'h0):(1'h0)])};
              reg132 <= reg128[(2'h2):(1'h0)];
              reg133 <= (($signed(reg133) >= (8'hb2)) ?
                  $signed({reg124,
                      $unsigned($signed(forvar116))}) : forvar119[(3'h5):(2'h3)]);
            end
        end
      reg134 <= reg127[(1'h0):(1'h0)];
    end
  assign wire135 = reg129[(4'he):(4'hc)];
  assign wire136 = reg117;
  assign wire137 = reg134;
  always
    @(posedge clk) begin
      reg138 <= $signed({(7'h41), reg115[(3'h4):(2'h3)]});
      if ((~^{reg127[(1'h0):(1'h0)], $unsigned((~&(wire113 > reg130)))}))
        begin
          for (forvar139 = (1'h0); (forvar139 < (2'h2)); forvar139 = (forvar139 + (1'h1)))
            begin
              reg140 <= wire114[(1'h0):(1'h0)];
            end
          if ($signed($unsigned({(reg123[(4'hf):(4'hc)] ?
                  wire112[(3'h4):(3'h4)] : {wire114}),
              reg140[(2'h3):(2'h2)]})))
            begin
              reg141 <= reg117[(1'h0):(1'h0)];
              reg142 = (-$signed($signed(reg132[(3'h4):(2'h3)])));
            end
          else
            begin
              reg141 <= reg141[(1'h1):(1'h0)];
              reg142 <= reg134[(2'h2):(1'h1)];
            end
          for (forvar143 = (1'h0); (forvar143 < (3'h4)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 <= ((8'hb4) >= wire110);
              reg145 <= wire136;
              reg146 = {$signed({"5Q2FWRsr7v",
                      $unsigned(reg118[(4'ha):(4'h8)])}),
                  reg124[(4'he):(4'hc)]};
              reg147 = $unsigned(reg118);
              reg148 <= $unsigned(reg120[(5'h10):(3'h4)]);
            end
        end
      else
        begin
          reg139 <= (reg127 ?
              $unsigned(wire113) : (($unsigned("cZfxgiVz0MM6yxn6Bs") ~^ (~^$signed((8'ha8)))) ?
                  reg126 : (8'h9d)));
          reg140 = (8'hb4);
        end
      for (forvar149 = (1'h0); (forvar149 < (3'h4)); forvar149 = (forvar149 + (1'h1)))
        begin
          reg150 <= ($unsigned($unsigned(reg121[(1'h1):(1'h0)])) ?
              (~&(~$unsigned($signed(reg131)))) : reg131[(4'h8):(3'h7)]);
        end
      if ((^~reg145[(3'h7):(2'h2)]))
        begin
          reg151 <= (8'hb1);
          for (forvar152 = (1'h0); (forvar152 < (1'h1)); forvar152 = (forvar152 + (1'h1)))
            begin
              reg153 = $unsigned(((8'hba) ? (8'hbd) : (~reg138)));
              reg154 <= {$unsigned(reg153[(2'h2):(2'h2)]), (~^(8'haf))};
              reg155 = "k8BzeF8L8rzLDTUM6";
              reg156 <= reg122;
            end
        end
      else
        begin
          reg151 <= ({(~{$unsigned(reg134)}),
              (forvar139 ?
                  reg139[(3'h4):(2'h3)] : $signed($signed(reg127)))} - (reg138[(4'hb):(3'h7)] <= ($signed(reg126) ?
              (8'hb0) : $signed(forvar149))));
          reg152 <= wire135[(3'h4):(2'h3)];
          for (forvar153 = (1'h0); (forvar153 < (2'h2)); forvar153 = (forvar153 + (1'h1)))
            begin
              reg154 <= $unsigned($signed((($signed(reg117) | {(8'hb8),
                  (8'hbb)}) <<< (&reg145))));
              reg155 <= (((($signed((7'h42)) ?
                          ((8'hae) >= (8'haa)) : forvar153) ^ reg124[(1'h1):(1'h1)]) ?
                      reg139 : (forvar152[(1'h1):(1'h0)] || $unsigned({(8'hb2)}))) ?
                  $signed($signed({(reg140 > (7'h41)),
                      (8'hb2)})) : (~reg147[(1'h0):(1'h0)]));
              reg156 <= (7'h43);
              reg157 <= forvar139;
            end
          for (forvar158 = (1'h0); (forvar158 < (2'h2)); forvar158 = (forvar158 + (1'h1)))
            begin
              reg159 <= reg118[(2'h3):(1'h1)];
              reg160 = {forvar119[(1'h0):(1'h0)]};
              reg161 <= $unsigned(forvar149);
              reg162 = reg133[(2'h3):(1'h1)];
              reg163 <= reg129;
            end
        end
      if (({((8'h9c) || (8'hb0)), (8'hbc)} != forvar149[(4'h8):(2'h3)]))
        begin
          reg164 <= (((reg161 && (~^reg123[(3'h5):(1'h0)])) >>> (((wire135 ?
                  wire111 : (8'hb3)) >>> $unsigned(reg152)) ?
              (!(8'hb9)) : $unsigned((reg141 ?
                  reg145 : (7'h41))))) < $signed((reg129[(3'h7):(3'h4)] ?
              reg159[(2'h3):(1'h0)] : reg154[(2'h2):(1'h0)])));
          reg165 <= {$unsigned($unsigned(forvar116[(1'h0):(1'h0)]))};
          reg166 = (((8'ha5) & ((^((8'hbe) || (8'hac))) + reg129)) == forvar153);
          reg167 = reg115[(1'h1):(1'h1)];
        end
      else
        begin
          for (forvar164 = (1'h0); (forvar164 < (2'h3)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 = reg163;
              reg166 <= ((8'hab) ^ forvar125[(5'h11):(4'hd)]);
            end
          if ($signed(forvar149))
            begin
              reg167 <= (((($unsigned((8'hae)) || $unsigned(reg150)) ?
                  (((8'h9d) < reg155) + (wire114 >>> reg138)) : ($unsigned(forvar116) ?
                      (reg152 | reg155) : $unsigned(reg130))) << reg159[(3'h6):(3'h5)]) >= forvar164[(4'ha):(3'h7)]);
            end
          else
            begin
              reg167 = $signed(reg121);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar168 = (1'h0); (forvar168 < (1'h0)); forvar168 = (forvar168 + (1'h1)))
        begin
          if ($unsigned(reg163))
            begin
              reg169 = forvar119;
              reg170 <= (({$unsigned((reg124 ? reg160 : (8'ha7)))} ?
                      ((forvar152 < {reg154,
                          (8'hab)}) == $unsigned((reg122 >> reg124))) : reg131[(3'h5):(2'h2)]) ?
                  wire136 : {forvar125, ((-reg167[(3'h5):(3'h5)]) << reg169)});
            end
          else
            begin
              reg169 <= ({{reg132}} < $unsigned(({{reg131, wire110},
                      reg161[(3'h6):(1'h0)]} ?
                  $unsigned($signed(reg118)) : {reg151, (8'hae)})));
              reg170 <= (reg169 - ((8'hb6) ?
                  reg142 : $unsigned(reg144[(5'h12):(3'h4)])));
              reg171 <= {{((8'hae) ^~ $unsigned($signed(forvar168)))},
                  (&(^~$unsigned({reg164})))};
              reg172 <= reg126;
              reg173 <= (~|reg150[(4'he):(2'h2)]);
            end
          if ($unsigned((^~(&(|forvar125[(3'h5):(3'h4)])))))
            begin
              reg174 = $signed($signed($signed((reg167 * (forvar164 ?
                  reg124 : (8'ha5))))));
              reg175 <= reg159[(2'h3):(2'h3)];
              reg176 = reg157;
              reg177 = reg121;
            end
          else
            begin
              reg174 <= (~&reg157);
              reg175 <= reg127;
              reg176 <= (reg151[(1'h0):(1'h0)] ~^ $signed(reg123[(4'hd):(4'hd)]));
              reg177 = (8'ha1);
              reg178 = {(((wire137 >> ((8'h9d) > forvar119)) + reg147[(1'h1):(1'h1)]) ?
                      (~|(wire111 || (forvar116 >>> wire136))) : (reg126 | {{(8'hac),
                              reg171}}))};
            end
          reg179 <= $unsigned(($signed((8'haf)) >>> (wire114[(2'h2):(1'h1)] * $signed((~reg171)))));
        end
      for (forvar180 = (1'h0); (forvar180 < (1'h0)); forvar180 = (forvar180 + (1'h1)))
        begin
          if ($unsigned(($signed((wire111[(4'hc):(2'h3)] ^ {reg144})) * (8'hb7))))
            begin
              reg181 <= $unsigned(reg179[(3'h7):(3'h6)]);
              reg182 <= $unsigned({(8'hac), (|reg163[(2'h2):(2'h2)])});
              reg183 <= reg167[(3'h4):(2'h2)];
              reg184 <= (reg146 <= reg172[(4'he):(3'h4)]);
            end
          else
            begin
              reg181 = $unsigned({{($unsigned(reg148) ?
                          (^(8'ha4)) : (8'hb0))}});
              reg182 <= reg184;
            end
        end
      for (forvar185 = (1'h0); (forvar185 < (1'h0)); forvar185 = (forvar185 + (1'h1)))
        begin
          reg186 <= {($unsigned(reg179) ?
                  $signed((((8'hb0) > reg147) ?
                      $signed((8'hb8)) : (forvar152 - reg147))) : reg154[(3'h4):(1'h1)])};
          if (reg167)
            begin
              reg187 <= reg169;
              reg188 = reg174;
            end
          else
            begin
              reg187 <= forvar139[(5'h13):(4'hf)];
              reg188 = reg183;
              reg189 <= {(reg175 ?
                      (reg150[(1'h0):(1'h0)] << $unsigned(reg173)) : (~^reg165))};
              reg190 = ({$unsigned(((~reg179) ?
                      $unsigned(forvar164) : {reg187})),
                  forvar149[(1'h1):(1'h1)]} << ((((|reg148) | {reg170,
                  reg129}) <= (reg117 ^ (|reg140))) + $unsigned(reg151)));
              reg191 <= reg151;
            end
        end
      reg192 <= {$unsigned($unsigned($signed({reg139, (8'hba)}))),
          ((reg146[(3'h4):(3'h4)] >>> {$signed((8'hbb))}) >> reg151)};
      for (forvar193 = (1'h0); (forvar193 < (3'h4)); forvar193 = (forvar193 + (1'h1)))
        begin
          reg194 = {(^~$signed({(forvar116 != reg128)})),
              $signed($signed(($unsigned(forvar139) << reg178[(3'h5):(3'h4)])))};
          if ($unsigned(((reg179 <= $unsigned(reg159)) ?
              {(|(reg182 ? reg152 : reg130)),
                  (^~((7'h42) ? reg152 : reg191))} : ("TYW" ?
                  reg123[(4'he):(4'hc)] : reg167[(1'h0):(1'h0)]))))
            begin
              reg195 = $unsigned($signed($unsigned(((!reg144) ?
                  (+forvar153) : reg148))));
              reg196 <= $unsigned((|(((forvar116 ?
                  reg175 : reg188) ^ forvar158[(4'h9):(1'h1)]) >= $signed("kVG3dVuMhyRAEQZp"))));
              reg197 <= {(8'hbe)};
              reg198 = reg174[(4'hb):(3'h6)];
            end
          else
            begin
              reg195 <= wire137;
              reg196 = reg192;
              reg197 = reg132;
              reg198 = "F1pFabmJ9R6w4MwU";
              reg199 <= ($signed(reg156) ?
                  (reg171[(4'ha):(3'h6)] ?
                      $unsigned({(reg161 ~^ forvar185),
                          (forvar125 ?
                              (8'hb1) : (8'hb5))}) : forvar139[(4'hd):(2'h3)]) : reg144);
            end
          for (forvar200 = (1'h0); (forvar200 < (1'h1)); forvar200 = (forvar200 + (1'h1)))
            begin
              reg201 <= ((8'ha2) >= ($signed($unsigned(((8'hb0) ^~ (8'hbd)))) <<< $unsigned({$signed(wire110),
                  forvar153})));
              reg202 <= ({(~&{(~^forvar168)})} ?
                  reg194 : {reg170[(4'hb):(4'ha)], reg188[(2'h2):(1'h0)]});
              reg203 <= "Yq7iCquk0nFtVC1M3opJ";
              reg204 <= reg178[(3'h6):(1'h1)];
            end
          for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
            begin
              reg206 = (8'hb0);
              reg207 <= reg203[(3'h5):(2'h3)];
              reg208 <= {((reg165[(3'h7):(2'h3)] * (reg144 << ((7'h42) + reg117))) ?
                      ((&(reg192 ?
                          reg202 : reg196)) * reg129) : {($unsigned(reg164) == {reg140,
                              (7'h40)}),
                          reg188}),
                  forvar152};
              reg209 <= reg182[(3'h4):(3'h4)];
            end
          for (forvar210 = (1'h0); (forvar210 < (2'h2)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= $unsigned($unsigned({(~^$signed((8'ha4))),
                  {{(8'hab), reg179}}}));
            end
        end
    end
  assign wire212 = (7'h44);
  always
    @(posedge clk) begin
      if (({reg195} != $unsigned($unsigned((-reg209[(1'h0):(1'h0)])))))
        begin
          reg213 = $unsigned((reg204[(2'h3):(1'h1)] ^ {($unsigned((8'ha5)) & $signed((8'hab))),
              reg173[(4'hc):(2'h2)]}));
          reg214 <= ((8'hba) > {(((reg183 << (8'ha9)) >= $unsigned((8'hb9))) ?
                  ((^reg139) >= (forvar152 <= reg183)) : "BGZ3")});
          reg215 <= forvar200;
          if (reg177)
            begin
              reg216 <= reg177[(4'ha):(4'h9)];
              reg217 <= ({$unsigned({reg181[(5'h13):(3'h6)], {reg121}}),
                  ({$unsigned(forvar143), ((8'hb9) ? (8'ha7) : (8'ha1))} ?
                      ($signed((8'hbf)) >= reg123) : $signed((reg166 < reg118)))} <= {$signed({reg201[(2'h2):(1'h0)]}),
                  reg146[(2'h2):(1'h0)]});
            end
          else
            begin
              reg216 <= $unsigned("NBybbIYhZzAyk");
              reg217 <= $signed(reg198[(1'h0):(1'h0)]);
              reg218 = (8'hae);
            end
        end
      else
        begin
          reg213 = $unsigned($unsigned(reg156[(4'h8):(3'h4)]));
          reg214 <= (reg138[(4'h9):(3'h6)] ^~ (^~{wire113}));
        end
      for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
        begin
          reg220 = (~&(+(8'hab)));
        end
      if ($unsigned(reg126[(2'h2):(1'h1)]))
        begin
          reg221 <= {{{(((8'hbd) > reg187) ?
                          {reg167} : reg134[(2'h3):(1'h1)])}}};
          reg222 <= reg187;
          reg223 = (~{(reg217 - forvar193[(2'h3):(1'h0)]),
              $unsigned({(reg192 >>> (7'h40))})});
          reg224 <= reg217;
          reg225 <= (reg128 ^ "l2HDEVdHIbeaB8eO");
        end
      else
        begin
          reg221 <= reg222;
          if ($unsigned({$unsigned(reg166)}))
            begin
              reg222 <= ($unsigned((($unsigned(forvar139) ?
                      (reg223 && reg132) : $signed((8'h9e))) + (8'hb5))) ?
                  $unsigned(reg194[(5'h10):(4'he)]) : $signed(($signed(reg216[(4'hc):(2'h2)]) ?
                      (8'ha8) : (~((8'ha1) ? (8'hbf) : (8'ha4))))));
            end
          else
            begin
              reg222 <= wire113;
              reg223 <= reg207[(1'h1):(1'h0)];
              reg224 = $unsigned(((~|(7'h43)) ?
                  reg166 : (reg175[(1'h0):(1'h0)] && (8'hbf))));
              reg225 = $signed($unsigned((&reg224[(1'h0):(1'h0)])));
              reg226 = (reg148 ?
                  {($unsigned((reg131 <= reg224)) ?
                          ((^forvar180) * (reg117 <<< reg225)) : (^~{reg140})),
                      (((7'h42) > ((8'haf) ?
                          (8'hba) : reg129)) ^~ {$signed(reg144)})} : $unsigned(forvar205[(4'ha):(1'h1)]));
            end
          reg227 <= (^~reg189);
        end
    end
  assign wire228 = {$signed(reg128[(2'h2):(1'h1)]),
                       {$unsigned({$signed(reg144)})}};
  assign wire229 = wire113;
  assign wire230 = $signed($unsigned((8'h9e)));
  assign wire231 = $signed(forvar210[(2'h3):(1'h0)]);
  always
    @(posedge clk) begin
      reg232 = {(({reg151, $unsigned(reg152)} * {$unsigned(reg148)}) ?
              ({$unsigned(reg142),
                  (8'hb4)} ^~ reg225[(2'h2):(1'h1)]) : "pKhzP")};
      reg233 = (forvar158[(4'hb):(3'h6)] != ($unsigned($signed({reg217,
          reg198})) | (-$unsigned(((8'ha3) ? reg218 : (8'h9e))))));
      if (reg224)
        begin
          for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 = (reg192 ?
                  (8'h9e) : (reg170 << {{(8'hb6), reg151[(3'h7):(2'h2)]}}));
            end
          reg236 = $signed(({{(~&reg151)}} < $unsigned(({reg221,
              (8'hbf)} ^~ wire230[(4'hb):(3'h6)]))));
          if ($unsigned(reg218))
            begin
              reg237 <= ({wire229[(1'h1):(1'h0)]} ^ reg218[(3'h5):(1'h1)]);
              reg238 <= ({(forvar125 ?
                          ("aLYpsbQ6zkYsng" <= reg165) : $signed((reg150 - reg157))),
                      (("I" || ((8'ha0) - reg222)) ^~ forvar158)} ?
                  reg201 : $unsigned($unsigned($unsigned({reg129,
                      forvar193}))));
              reg239 = reg179[(5'h13):(1'h1)];
            end
          else
            begin
              reg237 <= reg146[(4'ha):(1'h0)];
              reg238 <= forvar143;
              reg239 <= {(reg178[(3'h7):(1'h1)] || wire231),
                  {{$signed({forvar158, reg195}), reg182[(4'h9):(3'h5)]}}};
              reg240 <= ((8'ha4) >= $unsigned({((forvar219 ?
                      reg176 : reg238) ~^ (~|reg197))}));
            end
        end
      else
        begin
          reg234 = $signed((8'hbc));
          reg235 <= ((forvar234 && reg216) - $signed(forvar164[(3'h5):(3'h4)]));
          for (forvar236 = (1'h0); (forvar236 < (3'h4)); forvar236 = (forvar236 + (1'h1)))
            begin
              reg237 <= (7'h41);
              reg238 = $unsigned("G1thKiREMkVM");
            end
          for (forvar239 = (1'h0); (forvar239 < (2'h2)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= $unsigned("K");
              reg241 <= $unsigned($unsigned(forvar149[(1'h0):(1'h0)]));
              reg242 <= reg167;
            end
          for (forvar243 = (1'h0); (forvar243 < (2'h2)); forvar243 = (forvar243 + (1'h1)))
            begin
              reg244 <= {reg234,
                  ((forvar116 >= (^~$signed((8'haf)))) + (~|($signed(reg173) && $unsigned(reg141))))};
            end
        end
    end
  always
    @(posedge clk) begin
      reg245 <= (8'ha6);
      for (forvar246 = (1'h0); (forvar246 < (1'h0)); forvar246 = (forvar246 + (1'h1)))
        begin
          reg247 <= reg197;
        end
      for (forvar248 = (1'h0); (forvar248 < (1'h0)); forvar248 = (forvar248 + (1'h1)))
        begin
          for (forvar249 = (1'h0); (forvar249 < (2'h3)); forvar249 = (forvar249 + (1'h1)))
            begin
              reg250 = $unsigned(reg175);
              reg251 = "vMzOtdCdmJdL";
            end
          reg252 <= reg153[(1'h0):(1'h0)];
          for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= ($unsigned(reg201) == (-$signed((^reg142[(4'hc):(4'h8)]))));
              reg255 = forvar253[(2'h3):(2'h2)];
              reg256 = $unsigned($unsigned({((reg129 ? (8'hb6) : reg179) ?
                      (wire137 <<< reg244) : {reg250})}));
              reg257 <= (8'h9d);
              reg258 <= reg227[(2'h3):(2'h2)];
            end
        end
      reg259 <= ($unsigned(reg220[(4'hd):(1'h1)]) || ((((^forvar185) >= reg171[(4'hb):(3'h6)]) ?
          ((forvar246 ^ wire229) ?
              (reg254 <= forvar246) : (reg208 ?
                  (8'ha3) : (8'ha1))) : reg238[(1'h0):(1'h0)]) <= $signed((-reg154[(1'h0):(1'h0)]))));
    end
  assign wire260 = $signed((reg144[(2'h3):(1'h1)] ?
                       (($signed((8'h9d)) ?
                           $signed((8'hbb)) : $unsigned(reg177)) ~^ $signed({reg142})) : $signed((|reg215[(5'h10):(3'h4)]))));
  assign wire261 = (8'hb9);
  assign wire262 = $unsigned(reg178);
  assign wire263 = $unsigned((&$unsigned(((forvar180 < (8'hac)) - (^~reg134)))));
  assign wire264 = $signed($signed(((((8'ha5) >> forvar116) ?
                           (^~(8'hb7)) : (!reg138)) ?
                       ($signed(reg128) <<< reg204[(4'h8):(3'h5)]) : ($unsigned(reg255) | reg128))));
  assign wire265 = ({$unsigned(forvar205[(5'h13):(3'h4)])} ?
                       reg161[(4'ha):(1'h0)] : ((+$signed(((8'ha4) == reg227))) <= $signed(reg188)));
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param701 = (-(|((~|(^~(8'hb7))) ^ (((8'hac) ? (8'haa) : (8'h9d)) & (8'hbc)))))
, parameter param702 = (+{param701, {(-((8'h9c) >>> param701)), ((param701 ? (7'h43) : (8'h9f)) || (param701 << param701))}}) )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h6e3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire0;
  input wire [(5'h10):(1'h0)] wire1;
  input wire [(4'hc):(1'h0)] wire2;
  input wire signed [(5'h10):(1'h0)] wire3;
  reg signed [(4'ha):(1'h0)] reg700 = (1'h0);
  reg [(3'h4):(1'h0)] reg699 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg698 = (1'h0);
  reg [(3'h7):(1'h0)] reg697 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg696 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar695 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg694 = (1'h0);
  reg [(4'hd):(1'h0)] forvar693 = (1'h0);
  reg [(4'he):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg691 = (1'h0);
  reg [(4'ha):(1'h0)] reg690 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg689 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar688 = (1'h0);
  reg [(3'h7):(1'h0)] reg687 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar686 = (1'h0);
  reg [(4'he):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg684 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg683 = (1'h0);
  reg [(3'h7):(1'h0)] reg682 = (1'h0);
  reg [(4'h9):(1'h0)] reg681 = (1'h0);
  reg [(4'he):(1'h0)] reg680 = (1'h0);
  reg [(4'h8):(1'h0)] reg679 = (1'h0);
  reg [(4'hd):(1'h0)] reg678 = (1'h0);
  reg [(4'hf):(1'h0)] forvar677 = (1'h0);
  reg [(4'h9):(1'h0)] reg676 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire675;
  wire signed [(5'h11):(1'h0)] wire673;
  reg [(3'h4):(1'h0)] reg672 = (1'h0);
  reg [(4'hc):(1'h0)] reg671 = (1'h0);
  reg [(4'he):(1'h0)] reg670 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg669 = (1'h0);
  reg [(5'h13):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg666 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar665 = (1'h0);
  reg [(2'h2):(1'h0)] reg664 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg663 = (1'h0);
  reg [(5'h11):(1'h0)] reg662 = (1'h0);
  reg [(3'h4):(1'h0)] forvar661 = (1'h0);
  reg [(2'h2):(1'h0)] reg660 = (1'h0);
  reg [(4'hc):(1'h0)] reg659 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar658 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar657 = (1'h0);
  reg [(4'hd):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire5;
  wire signed [(4'hf):(1'h0)] wire6;
  wire [(5'h10):(1'h0)] wire553;
  reg signed [(4'ha):(1'h0)] forvar555 = (1'h0);
  reg [(4'hf):(1'h0)] reg556 = (1'h0);
  reg [(5'h12):(1'h0)] forvar557 = (1'h0);
  reg [(4'hc):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg559 = (1'h0);
  reg signed [(4'he):(1'h0)] reg557 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar560 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar561 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg562 = (1'h0);
  reg [(5'h13):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg565 = (1'h0);
  reg [(3'h5):(1'h0)] reg566 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar567 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg568 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg569 = (1'h0);
  reg signed [(4'he):(1'h0)] reg570 = (1'h0);
  reg [(5'h10):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg572 = (1'h0);
  reg [(4'hf):(1'h0)] reg573 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg574 = (1'h0);
  reg [(4'h8):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg577 = (1'h0);
  reg [(3'h4):(1'h0)] reg578 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire579;
  wire signed [(5'h13):(1'h0)] wire580;
  wire signed [(2'h2):(1'h0)] wire582;
  reg [(4'hd):(1'h0)] forvar583 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar584 = (1'h0);
  reg [(4'hd):(1'h0)] reg585 = (1'h0);
  reg [(4'h8):(1'h0)] reg586 = (1'h0);
  reg [(2'h3):(1'h0)] reg587 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg588 = (1'h0);
  reg [(4'h8):(1'h0)] forvar589 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg592 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg593 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar587 = (1'h0);
  reg [(4'he):(1'h0)] reg589 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg594 = (1'h0);
  reg [(3'h4):(1'h0)] reg595 = (1'h0);
  reg [(3'h7):(1'h0)] reg596 = (1'h0);
  wire [(2'h3):(1'h0)] wire597;
  wire signed [(3'h4):(1'h0)] wire598;
  reg signed [(5'h14):(1'h0)] forvar600 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar601 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(3'h6):(1'h0)] reg603 = (1'h0);
  reg [(5'h13):(1'h0)] forvar604 = (1'h0);
  reg [(2'h3):(1'h0)] forvar605 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg606 = (1'h0);
  reg [(4'he):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg608 = (1'h0);
  reg [(3'h7):(1'h0)] reg609 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar610 = (1'h0);
  reg [(5'h10):(1'h0)] reg611 = (1'h0);
  reg [(5'h15):(1'h0)] forvar612 = (1'h0);
  reg [(3'h6):(1'h0)] reg613 = (1'h0);
  reg [(5'h14):(1'h0)] reg614 = (1'h0);
  reg [(3'h4):(1'h0)] reg615 = (1'h0);
  reg [(5'h14):(1'h0)] reg616 = (1'h0);
  reg [(5'h13):(1'h0)] reg617 = (1'h0);
  reg [(5'h12):(1'h0)] reg618 = (1'h0);
  reg [(5'h10):(1'h0)] forvar619 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg620 = (1'h0);
  reg [(4'hf):(1'h0)] reg621 = (1'h0);
  reg [(2'h2):(1'h0)] forvar622 = (1'h0);
  reg [(5'h15):(1'h0)] forvar623 = (1'h0);
  reg [(4'ha):(1'h0)] reg624 = (1'h0);
  reg [(5'h13):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg626 = (1'h0);
  reg [(5'h11):(1'h0)] reg627 = (1'h0);
  reg [(5'h13):(1'h0)] reg628 = (1'h0);
  reg [(4'h9):(1'h0)] reg629 = (1'h0);
  reg [(3'h6):(1'h0)] reg630 = (1'h0);
  reg [(5'h11):(1'h0)] reg631 = (1'h0);
  reg [(5'h10):(1'h0)] forvar632 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg633 = (1'h0);
  reg [(2'h2):(1'h0)] reg634 = (1'h0);
  reg [(4'hf):(1'h0)] reg635 = (1'h0);
  reg [(5'h11):(1'h0)] reg636 = (1'h0);
  reg [(4'hb):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar638 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg639 = (1'h0);
  reg [(5'h15):(1'h0)] reg640 = (1'h0);
  reg [(5'h12):(1'h0)] reg641 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar643 = (1'h0);
  reg [(5'h14):(1'h0)] reg644 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg645 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg646 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg647 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg648 = (1'h0);
  reg [(2'h2):(1'h0)] reg649 = (1'h0);
  reg [(4'ha):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg651 = (1'h0);
  reg [(5'h14):(1'h0)] reg652 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar641 = (1'h0);
  reg signed [(4'he):(1'h0)] reg643 = (1'h0);
  wire [(5'h10):(1'h0)] wire654;
  assign y = {reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 forvar695,
                 reg694,
                 forvar693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 forvar688,
                 reg687,
                 forvar686,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 forvar677,
                 reg676,
                 wire675,
                 wire673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 forvar667,
                 reg666,
                 forvar665,
                 reg664,
                 reg663,
                 reg662,
                 forvar661,
                 reg660,
                 reg659,
                 forvar658,
                 forvar657,
                 reg656,
                 reg4,
                 wire5,
                 wire6,
                 wire553,
                 forvar555,
                 reg556,
                 forvar557,
                 reg558,
                 reg559,
                 reg557,
                 forvar560,
                 forvar561,
                 reg562,
                 reg563,
                 reg564,
                 reg565,
                 reg566,
                 forvar567,
                 reg568,
                 reg569,
                 reg570,
                 reg571,
                 reg572,
                 reg573,
                 reg574,
                 reg575,
                 reg576,
                 reg577,
                 reg578,
                 wire579,
                 wire580,
                 wire582,
                 forvar583,
                 forvar584,
                 reg585,
                 reg586,
                 reg587,
                 reg588,
                 forvar589,
                 reg590,
                 reg591,
                 reg592,
                 reg593,
                 forvar587,
                 reg589,
                 reg594,
                 reg595,
                 reg596,
                 wire597,
                 wire598,
                 forvar600,
                 forvar601,
                 reg602,
                 reg603,
                 forvar604,
                 forvar605,
                 reg606,
                 reg607,
                 reg608,
                 reg609,
                 forvar610,
                 reg611,
                 forvar612,
                 reg613,
                 reg614,
                 reg615,
                 reg616,
                 reg617,
                 reg618,
                 forvar619,
                 reg620,
                 reg621,
                 forvar622,
                 forvar623,
                 reg624,
                 reg625,
                 reg626,
                 reg627,
                 reg628,
                 reg629,
                 reg630,
                 reg631,
                 forvar632,
                 reg633,
                 reg634,
                 reg635,
                 reg636,
                 reg637,
                 forvar638,
                 reg639,
                 reg640,
                 reg641,
                 reg642,
                 forvar643,
                 reg644,
                 reg645,
                 reg646,
                 reg647,
                 reg648,
                 reg649,
                 reg650,
                 reg651,
                 reg652,
                 reg653,
                 forvar641,
                 reg643,
                 wire654,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 = $signed(((wire1[(3'h7):(3'h4)] ~^ $unsigned(wire3)) == wire2));
    end
  assign wire5 = wire2;
  assign wire6 = $unsigned(((({wire3} | (wire1 ? wire1 : (7'h43))) ?
                     wire3 : (((8'ha2) == wire3) & wire2[(4'h9):(3'h5)])) < $unsigned($unsigned((~wire2)))));
  module7 modinst554 (.clk(clk), .wire11(wire0), .wire10(wire3), .wire9(wire1), .y(wire553), .wire8(wire2));
  always
    @(posedge clk) begin
      if (wire3)
        begin
          for (forvar555 = (1'h0); (forvar555 < (1'h1)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 = ({$signed($signed((wire5 ? forvar555 : forvar555))),
                      (~&$signed($unsigned((8'hab))))} ?
                  wire1[(3'h4):(2'h2)] : wire3[(4'hc):(3'h7)]);
            end
          for (forvar557 = (1'h0); (forvar557 < (2'h2)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 = ($signed(reg556[(3'h4):(1'h0)]) & wire2[(4'hb):(4'h8)]);
              reg559 <= $signed($signed(wire553[(4'h9):(2'h3)]));
            end
        end
      else
        begin
          for (forvar555 = (1'h0); (forvar555 < (1'h1)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 <= "MC6";
              reg557 <= $signed((wire6[(1'h0):(1'h0)] ?
                  (~&wire553[(3'h5):(3'h4)]) : wire553[(4'hb):(1'h1)]));
              reg558 = $signed(wire6);
              reg559 <= {$signed((~reg4[(4'he):(4'hb)])),
                  ($signed($signed((&wire6))) ^ wire1)};
            end
        end
      for (forvar560 = (1'h0); (forvar560 < (2'h2)); forvar560 = (forvar560 + (1'h1)))
        begin
          for (forvar561 = (1'h0); (forvar561 < (1'h0)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 = {({({wire3} << (+forvar557))} ?
                      $signed(($unsigned(wire0) - (wire5 ?
                          (8'hb9) : (8'h9e)))) : ((wire1 != wire553) ?
                          $signed(wire6) : (~^wire1[(4'h8):(3'h6)])))};
              reg563 <= (&($signed($unsigned((~^reg562))) ?
                  $signed(((reg562 ?
                      (8'hb3) : forvar557) | $signed(wire2))) : ((^{(8'ha7)}) < ((&wire553) ?
                      ((8'h9f) * forvar561) : (~^reg562)))));
              reg564 = (reg558 ?
                  reg556[(1'h1):(1'h0)] : $signed(("n0enDM8" ?
                      reg556[(3'h7):(2'h3)] : $unsigned(reg556))));
              reg565 = ($signed((forvar555 ?
                      forvar557[(1'h0):(1'h0)] : (~&{(8'hb5), wire3}))) ?
                  $signed({$unsigned((wire5 & (8'ha9)))}) : (+wire5[(4'ha):(1'h1)]));
              reg566 = reg4;
            end
          for (forvar567 = (1'h0); (forvar567 < (2'h2)); forvar567 = (forvar567 + (1'h1)))
            begin
              reg568 = $unsigned((({$unsigned(wire0), (reg557 <= wire5)} ?
                  forvar555 : {(^wire3),
                      (wire3 ? reg564 : forvar557)}) + (^~{$signed(reg559)})));
            end
          reg569 = ($signed({(forvar561 && reg562)}) ?
              $signed(reg565) : $unsigned(($unsigned(forvar561[(4'hc):(4'hc)]) | (((8'h9d) ^~ forvar567) <<< (forvar557 ?
                  reg556 : reg556)))));
          if (($signed(wire0[(4'h8):(1'h0)]) < ($signed("47Cfshn2JFcYZC0xz") ?
              wire3 : (wire3 ?
                  (wire5[(4'hb):(3'h7)] ~^ $unsigned(reg4)) : wire5[(5'h10):(3'h7)]))))
            begin
              reg570 <= $signed(reg566[(2'h2):(1'h1)]);
              reg571 <= {($unsigned({$unsigned((8'hbd))}) ?
                      (~^(reg556 ?
                          {(8'hbd)} : (wire6 ? reg565 : forvar557))) : reg562),
                  (wire3[(3'h4):(1'h0)] ?
                      reg565[(5'h11):(3'h4)] : (~reg557[(2'h2):(1'h0)]))};
              reg572 = $signed(reg563[(4'h8):(3'h6)]);
              reg573 <= forvar567;
              reg574 = "Z8A";
            end
          else
            begin
              reg570 = {wire553, "I2Ki3l1x8W5"};
              reg571 = (reg558[(1'h0):(1'h0)] || ((($signed(reg573) <<< $signed(wire0)) ?
                  reg562[(4'he):(4'hc)] : ((~&reg565) <<< (reg572 ?
                      wire1 : (7'h44)))) && wire6[(2'h3):(1'h1)]));
            end
          if (($signed($signed($unsigned($signed(wire553)))) >> $signed({reg562[(4'h9):(2'h2)],
              ((^~reg563) ? (~|reg559) : $unsigned(reg574))})))
            begin
              reg575 <= {"4UFfmR"};
              reg576 <= $unsigned((((8'hb1) ?
                      (!(~&wire6)) : $unsigned(wire553[(2'h3):(2'h3)])) ?
                  $signed(((&wire5) > {reg569})) : $signed(({reg565, reg566} ?
                      $unsigned(reg570) : {reg571}))));
            end
          else
            begin
              reg575 = (forvar557 ? (|{$unsigned((-reg557))}) : reg4);
              reg576 <= "iuIvfiedN";
              reg577 <= forvar560[(2'h3):(1'h1)];
              reg578 = wire2[(2'h3):(1'h1)];
            end
        end
    end
  assign wire579 = $signed((((forvar567[(5'h10):(4'hd)] ?
                       {reg557, reg575} : (reg571 ?
                           reg570 : reg575)) + $unsigned((reg577 ?
                       forvar561 : (8'ha7)))) | (+"vDLPTYIIo9CbMb6")));
  module239 modinst581 (wire580, clk, reg557, reg577, reg556, forvar567);
  assign wire582 = (^(+{(-reg569), reg562[(4'he):(1'h0)]}));
  always
    @(posedge clk) begin
      for (forvar583 = (1'h0); (forvar583 < (3'h4)); forvar583 = (forvar583 + (1'h1)))
        begin
          for (forvar584 = (1'h0); (forvar584 < (2'h2)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 = (!(8'ha4));
              reg586 = $signed(((($signed(reg573) == (+reg568)) <= (|(8'hb0))) ?
                  $signed(((wire582 + reg575) ?
                      {reg585,
                          (8'ha8)} : $signed(wire3))) : (-(&$unsigned(wire580)))));
            end
        end
      if (reg585[(2'h3):(2'h3)])
        begin
          reg587 = $unsigned(reg576[(4'ha):(3'h7)]);
          reg588 <= forvar567[(3'h7):(1'h1)];
          for (forvar589 = (1'h0); (forvar589 < (2'h3)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 = reg4[(4'h8):(3'h5)];
              reg591 = $signed(reg570[(4'hc):(3'h4)]);
              reg592 <= "vVzdrv";
              reg593 = {((+$unsigned($unsigned((8'hb6)))) <<< (~((8'hb4) & reg568[(3'h5):(1'h1)]))),
                  {({((8'h9e) ? reg575 : forvar561),
                          (~(8'hae))} << forvar583[(1'h1):(1'h0)]),
                      (+($unsigned(reg576) - {(8'hb9)}))}};
            end
        end
      else
        begin
          for (forvar587 = (1'h0); (forvar587 < (3'h4)); forvar587 = (forvar587 + (1'h1)))
            begin
              reg588 <= $signed((^(~&reg575[(4'h8):(2'h3)])));
              reg589 <= ($signed(reg585) ?
                  reg575[(1'h0):(1'h0)] : (wire2 ?
                      (~&reg558) : $signed(reg593)));
              reg590 <= ($signed(forvar587[(1'h1):(1'h0)]) | (reg558 - reg585));
              reg591 = (((7'h42) ?
                      ($signed(reg569[(1'h1):(1'h0)]) <= $unsigned(reg4)) : $signed(reg593)) ?
                  reg566[(3'h5):(2'h3)] : (7'h41));
            end
          reg592 = (($unsigned($signed(reg576[(3'h5):(2'h2)])) > reg588) <<< ({reg569} ^~ ($unsigned((reg578 ?
                  (8'ha1) : reg562)) ?
              $signed((reg569 <= forvar560)) : forvar557[(1'h0):(1'h0)])));
        end
      reg594 <= ($unsigned(reg571) ?
          (-(^~$signed((~^reg575)))) : $signed(((8'hb7) ^ (~(reg4 < reg563)))));
      reg595 <= reg563[(3'h6):(1'h1)];
      reg596 <= reg566;
    end
  assign wire597 = $unsigned($unsigned($signed(reg591[(4'hd):(3'h6)])));
  module239 modinst599 (.clk(clk), .wire242(reg568), .wire243(wire3), .wire240(wire1), .y(wire598), .wire241(reg573));
  always
    @(posedge clk) begin
      for (forvar600 = (1'h0); (forvar600 < (2'h2)); forvar600 = (forvar600 + (1'h1)))
        begin
          for (forvar601 = (1'h0); (forvar601 < (2'h2)); forvar601 = (forvar601 + (1'h1)))
            begin
              reg602 = (~^(!$signed($signed((~|reg587)))));
            end
          reg603 = "8pxO0JOF";
        end
      for (forvar604 = (1'h0); (forvar604 < (2'h2)); forvar604 = (forvar604 + (1'h1)))
        begin
          for (forvar605 = (1'h0); (forvar605 < (2'h2)); forvar605 = (forvar605 + (1'h1)))
            begin
              reg606 = (~(($unsigned({forvar560, reg572}) ?
                  $signed(reg603) : reg558) << $unsigned(reg562)));
              reg607 = (reg602[(2'h2):(1'h0)] >= reg565[(2'h3):(1'h1)]);
              reg608 = reg586;
              reg609 <= $signed($unsigned((-reg574[(3'h4):(1'h1)])));
            end
          for (forvar610 = (1'h0); (forvar610 < (2'h2)); forvar610 = (forvar610 + (1'h1)))
            begin
              reg611 = ($unsigned((8'ha4)) != forvar567[(3'h4):(1'h0)]);
            end
          for (forvar612 = (1'h0); (forvar612 < (1'h1)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 <= reg578[(1'h0):(1'h0)];
              reg614 = $unsigned(wire597);
              reg615 <= $unsigned((reg563 * reg565[(5'h10):(3'h5)]));
              reg616 = $unsigned($signed((-reg558[(1'h0):(1'h0)])));
              reg617 = forvar601[(3'h5):(3'h5)];
            end
          reg618 = (8'hb1);
          for (forvar619 = (1'h0); (forvar619 < (3'h4)); forvar619 = (forvar619 + (1'h1)))
            begin
              reg620 = (({$signed((~|wire0))} ?
                      reg589 : ($signed(reg559) ?
                          $signed($unsigned(reg570)) : (!{forvar567}))) ?
                  wire2[(2'h2):(1'h1)] : reg578[(2'h3):(1'h1)]);
              reg621 <= $unsigned(((-reg559[(1'h1):(1'h0)]) >>> $unsigned(wire580)));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar622 = (1'h0); (forvar622 < (2'h3)); forvar622 = (forvar622 + (1'h1)))
        begin
          for (forvar623 = (1'h0); (forvar623 < (2'h2)); forvar623 = (forvar623 + (1'h1)))
            begin
              reg624 <= (8'hab);
              reg625 = $signed(reg558[(2'h2):(2'h2)]);
            end
          if ({(reg602 ?
                  (reg618[(4'he):(4'hd)] ?
                      (forvar623[(1'h1):(1'h1)] ?
                          (reg566 ?
                              wire1 : reg592) : $signed(reg591)) : $unsigned((reg4 << reg616))) : reg620[(3'h6):(3'h6)]),
              $signed($signed($signed("oi4m2OF")))})
            begin
              reg626 <= {(^($unsigned(wire3[(1'h0):(1'h0)]) ?
                      ((wire2 & reg606) ? {reg614} : reg573) : reg621))};
              reg627 = forvar589[(3'h5):(2'h3)];
            end
          else
            begin
              reg626 = reg572;
              reg627 = forvar589;
              reg628 = reg556;
              reg629 = reg625;
              reg630 = $signed(reg629[(2'h3):(1'h0)]);
            end
          reg631 <= (~&reg614[(4'hf):(3'h6)]);
          for (forvar632 = (1'h0); (forvar632 < (3'h4)); forvar632 = (forvar632 + (1'h1)))
            begin
              reg633 <= $unsigned((~reg559));
              reg634 <= $unsigned((-reg615[(2'h2):(2'h2)]));
              reg635 <= (forvar560 ~^ (^$unsigned(reg556)));
              reg636 = ({{"1QObHg2NGhW3h0DPgWDY", {$signed((7'h42))}},
                      reg566[(2'h3):(1'h1)]} ?
                  (reg634[(1'h0):(1'h0)] ?
                      (~|(~&(~^reg572))) : forvar612) : forvar567);
              reg637 <= reg593;
            end
          for (forvar638 = (1'h0); (forvar638 < (2'h3)); forvar638 = (forvar638 + (1'h1)))
            begin
              reg639 = (reg608[(3'h5):(2'h2)] - $signed($unsigned((reg608 && wire579[(2'h3):(2'h3)]))));
            end
        end
      reg640 = reg602[(1'h0):(1'h0)];
      if (reg563)
        begin
          reg641 = $unsigned({"2ZH53"});
          reg642 <= ($signed($unsigned((&(forvar632 <<< (8'ha3))))) * $unsigned((($unsigned(reg587) * $unsigned(reg557)) ^~ {reg590,
              {reg4, (8'ha8)}})));
          for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
            begin
              reg644 = reg574[(3'h5):(3'h4)];
              reg645 = (~^"UlLUUfzIdwhA5K5N1l8u");
              reg646 = reg570;
              reg647 <= (^reg565[(3'h4):(2'h3)]);
              reg648 = $unsigned($signed((^~($unsigned(reg566) >>> (!reg647)))));
            end
          if ((reg576 ?
              (&(^("4EFvuxruxBJL" <<< (reg618 ?
                  reg603 : forvar561)))) : {(~reg587),
                  $unsigned((~&(|wire6)))}))
            begin
              reg649 = $signed({reg564});
              reg650 = $unsigned(wire1);
              reg651 = ($unsigned({reg573,
                      $signed((reg577 ? reg562 : (8'hbc)))}) ?
                  $signed(reg594) : "ahDKFsHmLNK");
              reg652 = (((~((reg607 | (8'ha7)) ? {(8'ha5)} : {forvar612})) ?
                  ((|(forvar623 ?
                      reg589 : (8'hab))) < reg607[(1'h0):(1'h0)]) : ((7'h43) ?
                      reg566[(3'h4):(3'h4)] : $signed($unsigned(reg650)))) < ($signed("3vxbGW4g2xxuNV8") ?
                  reg617[(4'hd):(4'hb)] : (((reg629 ~^ (8'hab)) ~^ reg562[(3'h5):(2'h2)]) ?
                      reg621 : "")));
              reg653 <= "LANZIS";
            end
          else
            begin
              reg649 = reg596[(2'h3):(1'h0)];
            end
        end
      else
        begin
          for (forvar641 = (1'h0); (forvar641 < (2'h3)); forvar641 = (forvar641 + (1'h1)))
            begin
              reg642 = $unsigned(($unsigned((~&reg564)) ?
                  $unsigned(((reg566 > forvar601) ?
                      (reg634 ^~ forvar555) : $signed(reg609))) : (!(^~(reg565 - reg642)))));
              reg643 = $signed($unsigned($signed(((~reg578) || (^forvar612)))));
              reg644 <= $unsigned((~^(-forvar587[(3'h5):(3'h5)])));
            end
        end
    end
  module358 modinst655 (.wire363(reg588), .y(wire654), .wire362(reg646), .clk(clk), .wire361(reg576), .wire359(forvar557), .wire360(reg628));
  always
    @(posedge clk) begin
      reg656 = {$signed($unsigned((~reg616[(4'hb):(2'h3)])))};
      for (forvar657 = (1'h0); (forvar657 < (1'h0)); forvar657 = (forvar657 + (1'h1)))
        begin
          for (forvar658 = (1'h0); (forvar658 < (1'h0)); forvar658 = (forvar658 + (1'h1)))
            begin
              reg659 <= reg616;
              reg660 <= reg650;
            end
          for (forvar661 = (1'h0); (forvar661 < (2'h3)); forvar661 = (forvar661 + (1'h1)))
            begin
              reg662 <= forvar587[(3'h4):(3'h4)];
              reg663 = wire5[(2'h2):(2'h2)];
            end
          reg664 <= "uDauA";
        end
      for (forvar665 = (1'h0); (forvar665 < (1'h1)); forvar665 = (forvar665 + (1'h1)))
        begin
          reg666 <= $signed(((~|forvar661) ?
              $unsigned((reg566 ?
                  {reg611, reg649} : reg587)) : $unsigned($unsigned((reg572 ?
                  reg603 : forvar643)))));
          for (forvar667 = (1'h0); (forvar667 < (1'h1)); forvar667 = (forvar667 + (1'h1)))
            begin
              reg668 <= {{$unsigned($signed((wire2 - (8'hb5))))},
                  wire2[(3'h6):(1'h0)]};
              reg669 <= (($unsigned(((^~reg621) ?
                      (reg571 ? reg586 : forvar619) : {reg577, reg614})) ?
                  ((-(^~forvar657)) ?
                      reg571 : $signed(reg566)) : $unsigned((~&$unsigned(forvar605)))) + {{(((8'hbc) - forvar587) << (wire654 >>> forvar641)),
                      ((reg626 == reg668) || reg609)},
                  forvar638[(5'h14):(3'h6)]});
              reg670 = (((~&$signed($signed(reg614))) != ((+{(8'ha5),
                      (8'hbb)}) + (8'hb6))) ?
                  reg641[(2'h3):(2'h2)] : reg576);
              reg671 = wire0[(3'h6):(3'h5)];
              reg672 <= (reg630 >= $unsigned((forvar623[(2'h3):(1'h1)] ?
                  reg616[(5'h13):(3'h5)] : ($signed((7'h41)) ?
                      $unsigned(forvar641) : (-reg576)))));
            end
        end
    end
  module239 modinst674 (.wire243(reg670), .wire241(forvar610), .wire242(reg662), .wire240(forvar619), .y(wire673), .clk(clk));
  assign wire675 = reg585[(4'hb):(1'h0)];
  always
    @(posedge clk) begin
      reg676 <= reg627;
      for (forvar677 = (1'h0); (forvar677 < (2'h2)); forvar677 = (forvar677 + (1'h1)))
        begin
          if ({((~&{(reg591 ? (7'h44) : reg592)}) ?
                  ("0LZ7ulMy3Q" ? reg566 : (~(~|forvar604))) : (^~(~^(reg645 ?
                      reg574 : reg642)))),
              (|(|$signed((|reg585))))})
            begin
              reg678 = reg616;
              reg679 = $signed(({reg624[(4'ha):(4'h8)],
                      $signed({reg676, forvar612})} ?
                  $unsigned(({wire6} ?
                      (-wire598) : $unsigned(reg625))) : $unsigned((8'hbd))));
              reg680 = forvar667[(5'h12):(5'h10)];
            end
          else
            begin
              reg678 <= ((reg596[(1'h1):(1'h1)] ?
                  {(reg642[(2'h2):(2'h2)] ?
                          $unsigned(reg647) : {wire582,
                              reg566})} : $signed((8'hab))) ^ (^reg557[(4'hb):(3'h7)]));
              reg679 = ((8'haf) & (8'haa));
              reg680 <= (^$unsigned((forvar677 | $unsigned((wire6 ?
                  (8'ha4) : reg621)))));
              reg681 = $signed((+$signed({reg569[(3'h6):(3'h6)]})));
              reg682 = $signed((+$unsigned($signed(reg659[(4'h9):(2'h3)]))));
            end
          reg683 = ("AORJw0hctgzn" ? reg634 : reg628[(5'h12):(4'h9)]);
          reg684 <= (^~$unsigned($signed(("5SI4z0Rt" ?
              (&reg558) : $signed(forvar583)))));
        end
      reg685 = ({reg663, reg617} <= $unsigned(reg611[(3'h4):(3'h4)]));
      for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
        begin
          reg687 = reg603[(3'h5):(1'h0)];
          for (forvar688 = (1'h0); (forvar688 < (3'h4)); forvar688 = (forvar688 + (1'h1)))
            begin
              reg689 <= $unsigned((($unsigned(forvar612[(2'h2):(1'h1)]) - ((^~forvar583) - $signed(wire2))) ^~ reg587));
              reg690 <= ($unsigned($signed((|(&reg556)))) ?
                  ($unsigned(($unsigned(forvar589) ?
                          $unsigned((8'ha1)) : (reg591 < reg558))) ?
                      (~&{"n"}) : {(|reg558),
                          ($signed(reg621) <<< (!reg663))}) : reg651);
              reg691 <= (reg592 <<< reg687);
            end
          reg692 <= wire598;
          for (forvar693 = (1'h0); (forvar693 < (1'h0)); forvar693 = (forvar693 + (1'h1)))
            begin
              reg694 = (($unsigned((+reg595)) <= (({(8'ha3)} != reg672[(1'h1):(1'h1)]) ^~ ($unsigned(forvar623) + {reg630}))) ?
                  ((^~"FgMxdbLeRs39c2") ?
                      reg4[(5'h11):(3'h6)] : "4nApU95q8nfZ") : (((&((8'hb2) <<< reg590)) + reg647[(1'h1):(1'h0)]) * (~&$signed((reg603 ?
                      reg660 : wire654)))));
            end
          for (forvar695 = (1'h0); (forvar695 < (2'h3)); forvar695 = (forvar695 + (1'h1)))
            begin
              reg696 = (8'hab);
              reg697 <= (8'hae);
              reg698 <= forvar688[(1'h1):(1'h1)];
              reg699 = (!{(reg689 && (reg697 > (~&forvar583)))});
            end
        end
      reg700 = ($unsigned(forvar641) ?
          $signed($signed({reg595[(3'h4):(2'h2)],
              (^(8'ha9))})) : (((reg683[(1'h1):(1'h1)] ?
                  (&(7'h42)) : $signed(reg629)) << (~|(reg613 ?
                  reg635 : forvar632))) ?
              $unsigned({reg573[(4'hd):(4'hb)]}) : (8'hb9)));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7
#( parameter param551 = (((+(&((8'ha9) > (8'ha3)))) | (~((~^(8'ha9)) ? {(8'ha0), (8'haf)} : ((8'hbb) ? (8'h9c) : (8'hac))))) && (-((((8'ha6) ? (8'h9e) : (8'ha2)) ? ((8'hb1) != (8'hbd)) : ((8'hb0) ^ (8'ha8))) ? {((8'ha6) ? (8'hb6) : (8'hbc))} : (((8'haa) ~^ (8'hb3)) ? ((7'h40) != (8'ha5)) : ((8'ha3) < (8'hbb))))))
, parameter param552 = (((((param551 ? param551 : param551) <= (8'ha3)) != (param551 == {param551, param551})) ? {((param551 + param551) ? (~&param551) : (^param551))} : (~((param551 ? param551 : param551) ? (param551 ? param551 : param551) : (~param551)))) ? (8'hb4) : param551) )
(y, clk, wire11, wire10, wire9, wire8);
  output wire [(32'h814):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire11;
  input wire [(5'h10):(1'h0)] wire10;
  input wire [(4'h9):(1'h0)] wire9;
  input wire [(4'hc):(1'h0)] wire8;
  wire signed [(2'h3):(1'h0)] wire453;
  wire signed [(5'h10):(1'h0)] wire357;
  wire signed [(4'hf):(1'h0)] wire356;
  reg [(3'h7):(1'h0)] reg355 = (1'h0);
  reg [(4'ha):(1'h0)] reg354 = (1'h0);
  reg [(4'hb):(1'h0)] reg353 = (1'h0);
  reg [(4'h8):(1'h0)] reg352 = (1'h0);
  reg [(5'h11):(1'h0)] forvar351 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar350 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg347 = (1'h0);
  reg [(5'h11):(1'h0)] reg346 = (1'h0);
  reg [(5'h12):(1'h0)] reg345 = (1'h0);
  reg [(4'hc):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar343 = (1'h0);
  reg [(3'h4):(1'h0)] reg342 = (1'h0);
  reg [(4'hd):(1'h0)] forvar341 = (1'h0);
  reg [(4'ha):(1'h0)] reg340 = (1'h0);
  reg [(2'h3):(1'h0)] reg339 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg336 = (1'h0);
  reg [(2'h3):(1'h0)] forvar335 = (1'h0);
  reg [(4'hb):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg333 = (1'h0);
  reg [(5'h11):(1'h0)] reg332 = (1'h0);
  reg [(5'h15):(1'h0)] reg331 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar330 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg328 = (1'h0);
  reg [(2'h2):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar326 = (1'h0);
  reg [(4'hf):(1'h0)] reg325 = (1'h0);
  reg [(5'h11):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg323 = (1'h0);
  reg [(4'h8):(1'h0)] reg322 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg321 = (1'h0);
  reg [(4'hb):(1'h0)] forvar320 = (1'h0);
  reg [(3'h6):(1'h0)] reg319 = (1'h0);
  reg signed [(4'he):(1'h0)] reg318 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar317 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar315 = (1'h0);
  reg [(5'h13):(1'h0)] forvar314 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire235;
  reg signed [(4'h9):(1'h0)] reg43 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(4'hf):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg39 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar38 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar37 = (1'h0);
  reg [(4'hc):(1'h0)] reg36 = (1'h0);
  reg [(5'h10):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg34 = (1'h0);
  reg [(5'h12):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg32 = (1'h0);
  reg [(5'h10):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar27 = (1'h0);
  reg [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg25 = (1'h0);
  reg [(5'h13):(1'h0)] reg24 = (1'h0);
  reg [(4'h8):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar22 = (1'h0);
  reg [(4'hc):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg21 = (1'h0);
  reg [(3'h5):(1'h0)] forvar20 = (1'h0);
  reg [(5'h11):(1'h0)] reg19 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg18 = (1'h0);
  reg [(4'ha):(1'h0)] reg17 = (1'h0);
  reg [(5'h11):(1'h0)] reg16 = (1'h0);
  reg [(5'h15):(1'h0)] reg15 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg14 = (1'h0);
  reg [(3'h5):(1'h0)] reg13 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar12 = (1'h0);
  wire [(4'h8):(1'h0)] wire237;
  wire [(3'h6):(1'h0)] wire238;
  wire signed [(4'hd):(1'h0)] wire257;
  wire [(5'h13):(1'h0)] wire312;
  reg signed [(5'h14):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg456 = (1'h0);
  reg [(4'hc):(1'h0)] reg457 = (1'h0);
  reg [(4'ha):(1'h0)] reg458 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg459 = (1'h0);
  reg [(3'h7):(1'h0)] reg460 = (1'h0);
  reg [(3'h6):(1'h0)] reg461 = (1'h0);
  reg [(5'h15):(1'h0)] forvar459 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg463 = (1'h0);
  reg [(3'h6):(1'h0)] reg464 = (1'h0);
  reg [(5'h10):(1'h0)] reg465 = (1'h0);
  reg [(5'h12):(1'h0)] reg466 = (1'h0);
  reg [(4'hb):(1'h0)] reg467 = (1'h0);
  reg [(4'hd):(1'h0)] reg468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg469 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar470 = (1'h0);
  reg [(4'h9):(1'h0)] reg471 = (1'h0);
  reg [(2'h3):(1'h0)] forvar472 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg473 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg [(4'ha):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg476 = (1'h0);
  reg [(3'h6):(1'h0)] reg477 = (1'h0);
  reg [(3'h4):(1'h0)] reg478 = (1'h0);
  reg [(3'h7):(1'h0)] reg472 = (1'h0);
  reg [(3'h4):(1'h0)] forvar474 = (1'h0);
  reg [(5'h13):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar480 = (1'h0);
  reg [(2'h2):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg482 = (1'h0);
  reg [(4'hd):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg484 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar485 = (1'h0);
  reg [(3'h7):(1'h0)] reg486 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg487 = (1'h0);
  reg [(5'h15):(1'h0)] reg488 = (1'h0);
  reg [(3'h6):(1'h0)] reg489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg490 = (1'h0);
  reg [(3'h4):(1'h0)] reg491 = (1'h0);
  reg [(5'h10):(1'h0)] reg492 = (1'h0);
  reg [(3'h6):(1'h0)] reg493 = (1'h0);
  reg [(4'hd):(1'h0)] reg494 = (1'h0);
  wire [(2'h3):(1'h0)] wire495;
  wire [(4'hf):(1'h0)] wire496;
  reg [(2'h2):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar498 = (1'h0);
  reg [(4'h8):(1'h0)] reg499 = (1'h0);
  reg [(4'hf):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg501 = (1'h0);
  reg [(2'h3):(1'h0)] forvar502 = (1'h0);
  reg [(4'hd):(1'h0)] reg503 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar507 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg509 = (1'h0);
  reg [(2'h2):(1'h0)] reg510 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg511 = (1'h0);
  reg [(2'h3):(1'h0)] reg512 = (1'h0);
  reg [(4'hb):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg514 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire515;
  wire [(2'h2):(1'h0)] wire516;
  wire signed [(3'h6):(1'h0)] wire517;
  reg signed [(3'h5):(1'h0)] forvar518 = (1'h0);
  reg [(4'h8):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar521 = (1'h0);
  reg [(2'h2):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg523 = (1'h0);
  reg [(4'he):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg525 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar526 = (1'h0);
  reg [(2'h2):(1'h0)] reg527 = (1'h0);
  reg [(3'h5):(1'h0)] reg528 = (1'h0);
  reg [(4'h9):(1'h0)] forvar529 = (1'h0);
  reg [(2'h2):(1'h0)] reg530 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg531 = (1'h0);
  reg [(5'h12):(1'h0)] forvar532 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg534 = (1'h0);
  reg [(4'hc):(1'h0)] forvar535 = (1'h0);
  reg [(5'h11):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg537 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg539 = (1'h0);
  reg [(4'hb):(1'h0)] forvar540 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg541 = (1'h0);
  reg [(4'hc):(1'h0)] reg542 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg544 = (1'h0);
  reg [(5'h14):(1'h0)] reg545 = (1'h0);
  reg [(5'h14):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg532 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg540 = (1'h0);
  reg [(2'h3):(1'h0)] reg547 = (1'h0);
  reg [(4'hd):(1'h0)] reg548 = (1'h0);
  wire [(2'h2):(1'h0)] wire549;
  assign y = {wire453,
                 wire357,
                 wire356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 forvar351,
                 forvar350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 forvar343,
                 reg342,
                 forvar341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 forvar335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 forvar330,
                 reg329,
                 reg328,
                 reg327,
                 forvar326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 forvar317,
                 reg316,
                 forvar315,
                 forvar314,
                 wire235,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 forvar38,
                 forvar37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 forvar27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 forvar22,
                 reg22,
                 reg21,
                 forvar20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 forvar12,
                 wire237,
                 wire238,
                 wire257,
                 wire312,
                 reg455,
                 reg456,
                 reg457,
                 reg458,
                 reg459,
                 reg460,
                 reg461,
                 forvar459,
                 reg462,
                 reg463,
                 reg464,
                 reg465,
                 reg466,
                 reg467,
                 reg468,
                 reg469,
                 forvar470,
                 reg471,
                 forvar472,
                 reg473,
                 reg474,
                 reg475,
                 reg476,
                 reg477,
                 reg478,
                 reg472,
                 forvar474,
                 reg479,
                 forvar480,
                 reg481,
                 reg482,
                 reg483,
                 reg484,
                 forvar485,
                 reg486,
                 reg487,
                 reg488,
                 reg489,
                 reg490,
                 reg491,
                 reg492,
                 reg493,
                 reg494,
                 wire495,
                 wire496,
                 reg497,
                 forvar498,
                 reg499,
                 reg500,
                 reg501,
                 forvar502,
                 reg503,
                 reg504,
                 reg505,
                 reg506,
                 forvar507,
                 reg508,
                 reg509,
                 reg510,
                 reg511,
                 reg512,
                 reg513,
                 reg514,
                 wire515,
                 wire516,
                 wire517,
                 forvar518,
                 reg519,
                 reg520,
                 forvar521,
                 reg522,
                 reg523,
                 reg524,
                 reg525,
                 forvar526,
                 reg527,
                 reg528,
                 forvar529,
                 reg530,
                 reg531,
                 forvar532,
                 reg533,
                 reg534,
                 forvar535,
                 reg536,
                 reg537,
                 reg538,
                 reg539,
                 forvar540,
                 reg541,
                 reg542,
                 reg543,
                 reg544,
                 reg545,
                 reg546,
                 reg532,
                 reg535,
                 reg540,
                 reg547,
                 reg548,
                 wire549,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar12 = (1'h0); (forvar12 < (1'h0)); forvar12 = (forvar12 + (1'h1)))
        begin
          if (($signed((forvar12 >>> ({forvar12} ?
                  ((8'haa) | wire10) : {wire9}))) ?
              (wire8[(3'h4):(1'h0)] ?
                  $signed(wire9[(2'h3):(1'h1)]) : wire9[(3'h6):(1'h1)]) : $signed(((-(!wire11)) ?
                  (^(wire8 ? wire9 : wire10)) : {(wire8 ? wire8 : forvar12)}))))
            begin
              reg13 <= $unsigned({(((wire8 - wire9) <<< wire10) ^~ ({wire11,
                          wire8} ?
                      wire10[(1'h1):(1'h1)] : (wire11 > (8'had)))),
                  ($signed((wire10 ? wire9 : wire11)) >= wire10)});
              reg14 <= $signed(wire10);
              reg15 = {reg13[(2'h3):(2'h3)], $unsigned((|(7'h42)))};
            end
          else
            begin
              reg13 <= wire8[(4'hc):(2'h2)];
              reg14 <= (|$unsigned((~&($unsigned(wire8) ? wire11 : reg14))));
              reg15 = {$unsigned(($signed(reg13) * ($unsigned((8'hbb)) ?
                      reg13[(2'h2):(1'h1)] : $signed(wire9)))),
                  $unsigned((~^"03iE0U"))};
              reg16 = $unsigned(wire9[(2'h3):(2'h3)]);
              reg17 <= {(&$unsigned($signed((reg13 * reg16))))};
            end
          reg18 = wire8[(4'h9):(2'h2)];
        end
      reg19 <= $signed(($signed($unsigned({forvar12, reg18})) ?
          (+(!reg17[(3'h4):(1'h0)])) : ((forvar12[(1'h0):(1'h0)] != ((8'hba) ?
                  forvar12 : reg15)) ?
              $unsigned(reg14) : $unsigned(((8'hbb) ~^ reg17)))));
      for (forvar20 = (1'h0); (forvar20 < (1'h0)); forvar20 = (forvar20 + (1'h1)))
        begin
          reg21 = forvar12;
        end
      if (forvar20)
        begin
          reg22 = reg17[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar22 = (1'h0); (forvar22 < (1'h0)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= $unsigned(($signed(((reg21 >= reg13) ?
                      forvar12[(1'h1):(1'h0)] : ((8'hbd) ? reg22 : wire8))) ?
                  ($unsigned({wire11, reg17}) ?
                      $unsigned(((8'hbf) ?
                          reg16 : (8'ha4))) : reg17[(2'h3):(2'h3)]) : reg22[(4'h8):(3'h5)]));
            end
          if ((forvar22 ^~ $signed(reg17[(2'h3):(2'h2)])))
            begin
              reg24 <= ((~|((|reg15[(3'h4):(3'h4)]) ?
                  wire10 : $unsigned((|reg13)))) <<< $signed((reg17[(1'h1):(1'h1)] ?
                  $unsigned(((7'h40) ? forvar22 : (8'ha4))) : reg16)));
              reg25 = (reg17 ?
                  {("1" ?
                          (&(reg21 > wire9)) : ((!(8'h9c)) ?
                              $signed((8'hb6)) : {wire10})),
                      ((forvar22 || $unsigned(forvar22)) ?
                          forvar20[(2'h3):(2'h3)] : $unsigned(reg17))} : $signed($unsigned({(&forvar12),
                      (~wire11)})));
              reg26 = (~&(!({(reg24 ? reg17 : (8'ha0))} ?
                  (^$signed((8'ha7))) : ((wire8 ? reg17 : reg18) < (reg14 ?
                      reg25 : wire10)))));
            end
          else
            begin
              reg24 = $unsigned($unsigned(reg19));
            end
          for (forvar27 = (1'h0); (forvar27 < (3'h4)); forvar27 = (forvar27 + (1'h1)))
            begin
              reg28 = {reg17, (&((|(~wire11)) ? reg13 : "y1DJpXmVEfV1qebQ"))};
              reg29 = $unsigned($signed((reg25[(1'h0):(1'h0)] <= wire9[(3'h5):(3'h4)])));
              reg30 <= $signed(reg29);
              reg31 <= reg19[(3'h6):(1'h0)];
            end
          reg32 = ($signed((~^{$unsigned((8'hac)),
              (reg16 ? reg29 : reg23)})) ~^ (&reg21));
          if (reg14)
            begin
              reg33 = (8'ha8);
              reg34 <= (8'h9c);
            end
          else
            begin
              reg33 = reg21;
              reg34 <= ($unsigned({(^((8'hb4) | (7'h41))),
                  $unsigned({forvar22})}) || (~|reg13));
              reg35 = (~|(wire10 <= (~^$unsigned((reg18 >> reg34)))));
              reg36 = reg19;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar37 = (1'h0); (forvar37 < (1'h1)); forvar37 = (forvar37 + (1'h1)))
        begin
          for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= $unsigned($signed($unsigned($unsigned($signed(reg14)))));
            end
          reg40 <= $unsigned(forvar37[(3'h7):(3'h6)]);
          reg41 = $signed(reg16[(4'h8):(2'h3)]);
        end
      if (reg19)
        begin
          reg42 <= (|$unsigned((8'h9c)));
          reg43 = (7'h44);
        end
      else
        begin
          reg42 = (+$unsigned($signed($signed(forvar37[(3'h7):(1'h0)]))));
        end
    end
  module44 modinst236 (wire235, clk, reg17, wire11, forvar37, reg33, reg16);
  assign wire237 = (&$signed($signed((reg18[(4'h9):(3'h4)] ?
                       ((8'hb3) ? reg29 : (8'haf)) : {wire235, forvar22}))));
  assign wire238 = reg26;
  module239 modinst258 (wire257, clk, reg34, reg24, forvar27, wire10);
  module259 modinst313 (.wire260(reg15), .clk(clk), .wire261(wire257), .y(wire312), .wire262(reg22), .wire263(reg34), .wire264(reg26));
  always
    @(posedge clk) begin
      for (forvar314 = (1'h0); (forvar314 < (1'h1)); forvar314 = (forvar314 + (1'h1)))
        begin
          for (forvar315 = (1'h0); (forvar315 < (3'h4)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 = $signed(((~&$unsigned((^reg22))) && $unsigned(wire257)));
            end
          for (forvar317 = (1'h0); (forvar317 < (2'h3)); forvar317 = (forvar317 + (1'h1)))
            begin
              reg318 = $unsigned($signed($unsigned($unsigned($unsigned((8'hac))))));
              reg319 = ($signed(reg21) >>> (($unsigned({forvar12}) <= ((reg17 ?
                  reg42 : wire237) <<< ((7'h41) ?
                  reg32 : (8'hbc)))) >>> (!reg13[(2'h3):(2'h3)])));
            end
          for (forvar320 = (1'h0); (forvar320 < (1'h1)); forvar320 = (forvar320 + (1'h1)))
            begin
              reg321 = $unsigned(reg42);
              reg322 = {(forvar38[(1'h1):(1'h1)] < reg18)};
              reg323 <= $signed($signed((reg22 ? reg25 : (~^reg14))));
              reg324 = $unsigned($signed($signed($unsigned(reg34[(4'h8):(3'h6)]))));
              reg325 <= (wire10[(4'hd):(4'hd)] == reg30);
            end
          for (forvar326 = (1'h0); (forvar326 < (1'h1)); forvar326 = (forvar326 + (1'h1)))
            begin
              reg327 = (|((^~forvar37) <= $signed($signed(reg318[(4'hd):(2'h2)]))));
              reg328 <= reg24[(5'h13):(3'h4)];
              reg329 <= forvar314[(4'h8):(3'h5)];
            end
        end
      for (forvar330 = (1'h0); (forvar330 < (2'h2)); forvar330 = (forvar330 + (1'h1)))
        begin
          if ($signed($unsigned(($unsigned((reg21 ?
              reg42 : forvar315)) - ($unsigned(reg13) ?
              (&reg325) : (-forvar20))))))
            begin
              reg331 <= wire10;
              reg332 = $unsigned((^(8'hb2)));
              reg333 <= ($signed((reg35 | "Yd")) ?
                  "cWWWhSJ53qD9SZsz6bKT" : reg19[(4'hc):(4'ha)]);
              reg334 <= {{reg325}};
            end
          else
            begin
              reg331 = $signed(wire8);
              reg332 <= $signed(reg323[(1'h1):(1'h1)]);
            end
          for (forvar335 = (1'h0); (forvar335 < (3'h4)); forvar335 = (forvar335 + (1'h1)))
            begin
              reg336 <= (((forvar326 ?
                      ((&wire238) ?
                          {reg331} : {reg29, (8'hac)}) : wire8[(3'h4):(1'h1)]) ?
                  (~$signed(forvar320[(1'h1):(1'h1)])) : (^~$unsigned(forvar330))) ~^ $signed($signed(forvar335)));
              reg337 = $unsigned($unsigned(reg319[(2'h3):(2'h3)]));
              reg338 <= forvar320;
              reg339 <= {reg329,
                  ((-$signed($signed(reg327))) ?
                      forvar314 : {((reg327 - (8'hb5)) ? "DaC1UJ" : (|reg31)),
                          (|(reg318 > reg319))})};
              reg340 <= {($unsigned($signed($signed(reg41))) ?
                      ({"pZICGkgBa"} ^~ $signed(((8'ha7) ?
                          (8'ha8) : reg329))) : (8'hb2))};
            end
          for (forvar341 = (1'h0); (forvar341 < (3'h4)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 = $signed(("2nJeSbMB9P" ?
                  reg40 : $unsigned($signed(reg332))));
            end
          for (forvar343 = (1'h0); (forvar343 < (1'h1)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 = $unsigned({$unsigned(reg21), reg338});
              reg345 = ($signed(((^~(&(7'h41))) ?
                  ((reg41 ? reg324 : reg14) ?
                      (reg333 ?
                          wire312 : reg336) : reg19) : (&reg340[(1'h0):(1'h0)]))) * (|reg332));
              reg346 = reg332;
            end
        end
      reg347 <= $unsigned({$signed(reg32)});
      reg348 = ({(!(((7'h40) <= reg324) || $signed((8'ha3)))),
          {((wire10 & wire10) & $unsigned(reg29))}} >> forvar315);
      reg349 = {{forvar317}};
    end
  always
    @(posedge clk) begin
      for (forvar350 = (1'h0); (forvar350 < (1'h0)); forvar350 = (forvar350 + (1'h1)))
        begin
          for (forvar351 = (1'h0); (forvar351 < (1'h0)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 = ($unsigned((((reg325 & reg340) >> forvar326[(5'h11):(4'hf)]) || reg331[(1'h1):(1'h1)])) ?
                  $unsigned(reg348[(3'h6):(2'h3)]) : (({{reg29}} ?
                          $signed($unsigned(forvar315)) : forvar38[(3'h4):(3'h4)]) ?
                      forvar326[(3'h5):(3'h4)] : $unsigned($signed((8'ha5)))));
              reg353 = ({(wire8 == wire238[(3'h4):(2'h2)]),
                  $unsigned($signed((reg327 ?
                      reg324 : forvar37)))} | (~&(reg21 | (!(~|reg39)))));
            end
        end
      reg354 = $signed(wire238);
      reg355 <= $signed($unsigned(($unsigned(reg32[(3'h4):(2'h3)]) << reg36[(1'h1):(1'h1)])));
    end
  assign wire356 = $signed($signed($signed(((forvar326 - reg333) ?
                       $signed(reg31) : reg334[(3'h5):(2'h3)]))));
  assign wire357 = {reg42[(1'h0):(1'h0)]};
  module358 modinst454 (wire453, clk, reg321, wire356, reg346, forvar315, wire312);
  always
    @(posedge clk) begin
      reg455 <= reg25;
      if (forvar335)
        begin
          if ($signed(reg16[(4'h8):(1'h1)]))
            begin
              reg456 = (~&(~|$unsigned(wire312)));
              reg457 <= (|(reg319 ?
                  reg324[(4'hf):(4'hf)] : $signed((~|(~wire10)))));
              reg458 = ($unsigned($signed(((|wire238) ^~ $signed(wire8)))) == ((($unsigned(reg456) >>> $unsigned(reg327)) ?
                      $unsigned((~&reg336)) : ($unsigned(reg345) ?
                          (+forvar12) : $unsigned(reg40))) ?
                  (((reg13 + reg348) <<< {reg29,
                      reg32}) << (^"DWNWrtzAFilRgT")) : (reg40 >>> reg42[(3'h4):(1'h1)])));
              reg459 = $signed((reg345[(3'h7):(1'h0)] << (|reg41[(3'h6):(2'h2)])));
              reg460 = ((+({(|wire357)} && reg23)) == (reg25 >= (8'had)));
            end
          else
            begin
              reg456 = (+$signed((($signed(forvar326) ?
                  (~&wire10) : $signed(reg33)) >> $signed((8'hb2)))));
            end
          reg461 = (reg319 ?
              wire11 : ($unsigned($signed(forvar326[(4'hf):(4'hf)])) ?
                  (^~(reg459[(1'h1):(1'h0)] ?
                      (forvar335 | reg329) : {(8'h9c),
                          reg354})) : ((|$signed((8'ha1))) >= $signed(((8'haf) >= reg322)))));
        end
      else
        begin
          reg456 = $signed(((8'ha2) | "4z6hJXctrTEHSGO"));
          reg457 <= (&$unsigned((~|((^wire356) ~^ reg33[(4'h8):(3'h7)]))));
          reg458 <= (+forvar38[(2'h3):(1'h0)]);
          for (forvar459 = (1'h0); (forvar459 < (2'h2)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 <= (-(^(~|($unsigned(wire10) >> (forvar330 & forvar20)))));
              reg461 <= reg318;
              reg462 = $signed((~|wire453[(1'h0):(1'h0)]));
              reg463 = (-($unsigned($signed({forvar37,
                  reg355})) - (wire235[(4'hf):(3'h5)] && reg333)));
              reg464 <= $unsigned((forvar317 ?
                  $signed({(reg347 >>> reg318)}) : $signed(reg21[(5'h10):(5'h10)])));
            end
          if ($signed(reg26[(4'hf):(3'h7)]))
            begin
              reg465 <= $signed({$unsigned((reg15[(3'h5):(3'h5)] ?
                      reg14[(2'h3):(1'h1)] : reg13))});
              reg466 <= $signed($signed((forvar27 || ($signed(reg21) ?
                  (forvar351 ? reg337 : reg322) : $signed(reg354)))));
            end
          else
            begin
              reg465 <= ((((&reg333) ^ ((^~reg23) >= $signed(forvar37))) >= wire237) ?
                  ((|$unsigned((forvar351 <= reg316))) ?
                      $signed((~forvar335[(2'h2):(2'h2)])) : (+($unsigned(reg461) && (-(8'hb7))))) : reg462[(1'h0):(1'h0)]);
              reg466 <= forvar314;
              reg467 <= reg322[(2'h2):(2'h2)];
              reg468 <= (((-(&((8'hbc) ? reg33 : reg460))) ?
                      $unsigned((wire312 != (&(8'h9d)))) : ($signed($signed(reg349)) ?
                          ($signed(reg33) != (~|forvar317)) : {(reg17 ?
                                  reg318 : reg336),
                              (^~reg43)})) ?
                  (($signed(((8'hb3) ? reg339 : (8'had))) ?
                          (forvar330[(2'h3):(2'h2)] ^ (wire356 <= reg325)) : reg353[(1'h0):(1'h0)]) ?
                      (((reg342 ? reg31 : wire8) ?
                              $signed(reg333) : $signed(forvar326)) ?
                          $signed((~|reg459)) : $unsigned($signed(reg13))) : (((reg329 || wire9) <<< forvar320[(3'h6):(1'h0)]) >= $unsigned($unsigned(wire356)))) : (!$unsigned(reg462)));
              reg469 <= "C";
            end
        end
      if ($unsigned(reg336[(3'h4):(3'h4)]))
        begin
          for (forvar470 = (1'h0); (forvar470 < (2'h2)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 <= $signed(($signed((8'ha4)) ?
                  {(wire8[(3'h6):(1'h1)] < "8s0ndD2kvTIxGSU38q"),
                      ("Cd4ZZv6SlctX" & forvar351[(3'h6):(1'h1)])} : $unsigned(reg333)));
            end
          for (forvar472 = (1'h0); (forvar472 < (1'h1)); forvar472 = (forvar472 + (1'h1)))
            begin
              reg473 <= $signed(reg325);
              reg474 = {$signed($unsigned(($signed(reg461) >>> (reg318 - forvar330)))),
                  reg14[(3'h4):(3'h4)]};
              reg475 <= (~{(^(reg344 + $unsigned(reg322))),
                  $signed(($unsigned(reg18) > (8'ha8)))});
              reg476 <= {reg354};
              reg477 <= ((+{{(forvar350 >>> reg473)},
                      $unsigned((reg457 ? reg464 : reg318))}) ?
                  $unsigned(reg468) : {(^((|reg22) != {(8'hbc), reg456}))});
            end
          reg478 = reg327[(1'h1):(1'h1)];
        end
      else
        begin
          for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 = forvar317[(2'h3):(2'h2)];
              reg472 <= reg476;
              reg473 = wire356;
            end
          for (forvar474 = (1'h0); (forvar474 < (1'h0)); forvar474 = (forvar474 + (1'h1)))
            begin
              reg475 = (reg340 - ($signed("wNORN6MgEJwOEzm") >>> reg34));
              reg476 <= $unsigned($unsigned($unsigned(forvar38)));
              reg477 = ($unsigned(forvar470) ? reg471[(2'h3):(2'h3)] : "BiR");
              reg478 = "8JQaVpWEtSRkZv";
              reg479 = $signed({$unsigned(((8'h9c) ?
                      (reg327 << reg458) : reg29[(1'h0):(1'h0)])),
                  reg15});
            end
          for (forvar480 = (1'h0); (forvar480 < (2'h2)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 = "Tp9";
              reg482 = (forvar341[(1'h1):(1'h1)] ?
                  $signed($unsigned($unsigned($unsigned(reg476)))) : reg462);
            end
          reg483 <= {($unsigned(reg33[(4'hd):(4'ha)]) & reg349[(1'h0):(1'h0)]),
              $unsigned($signed((!(reg21 ? forvar314 : reg466))))};
        end
      reg484 <= ($unsigned($signed(reg43)) ?
          (^~($unsigned(reg324[(5'h10):(4'hb)]) ?
              $signed($signed(reg469)) : $unsigned($signed(reg35)))) : $unsigned(reg347));
      for (forvar485 = (1'h0); (forvar485 < (2'h2)); forvar485 = (forvar485 + (1'h1)))
        begin
          if ($signed($unsigned(reg465[(4'ha):(2'h2)])))
            begin
              reg486 <= {({$signed((~&reg345)),
                      $signed($signed((8'ha3)))} | (reg471[(2'h2):(1'h0)] + $unsigned("Sr3R5w4Y")))};
              reg487 = ($unsigned((~&{(reg331 ? reg33 : reg462),
                  (-reg19)})) >> ((7'h42) ?
                  (~|$unsigned((~^(8'hae)))) : {$signed((+wire235)),
                      reg323[(1'h1):(1'h0)]}));
            end
          else
            begin
              reg486 <= (8'ha7);
              reg487 <= forvar472;
              reg488 <= $signed(reg465[(3'h6):(3'h5)]);
              reg489 <= wire237[(1'h1):(1'h0)];
            end
          reg490 <= {$unsigned(reg457),
              ($signed(forvar326) != (~$signed($unsigned(reg461))))};
          reg491 <= reg333[(4'ha):(4'h9)];
          if ((forvar343 ?
              ($signed(($unsigned(forvar470) ?
                      (reg465 ? reg31 : reg459) : reg328[(3'h6):(2'h2)])) ?
                  (+(~^((8'hac) ^~ reg34))) : $signed(($signed(forvar12) | (8'hb3)))) : (reg22 ~^ reg14[(1'h0):(1'h0)])))
            begin
              reg492 <= (reg461 ^~ $signed(reg39[(2'h3):(1'h0)]));
              reg493 <= {$unsigned((forvar12 ^~ $unsigned($signed(reg342)))),
                  $unsigned(forvar351[(2'h2):(1'h0)])};
              reg494 <= (8'ha4);
            end
          else
            begin
              reg492 = ($signed((&{$unsigned(reg458), forvar37})) ?
                  $signed($unsigned(((forvar470 != reg457) + $unsigned(reg489)))) : ($signed((|reg489)) ?
                      reg329[(3'h5):(3'h4)] : $signed($unsigned(reg29[(3'h7):(3'h6)]))));
              reg493 <= reg36;
            end
        end
    end
  assign wire495 = (7'h43);
  assign wire496 = {reg333,
                       ($unsigned(reg490[(4'h8):(1'h1)]) ^~ $unsigned({{reg329,
                               forvar317},
                           (reg348 ~^ reg32)}))};
  always
    @(posedge clk) begin
      reg497 <= reg33[(4'hb):(1'h0)];
      for (forvar498 = (1'h0); (forvar498 < (1'h0)); forvar498 = (forvar498 + (1'h1)))
        begin
          if ($unsigned($signed($unsigned($unsigned(reg353)))))
            begin
              reg499 <= ($unsigned((($signed(wire237) ?
                  $unsigned(reg483) : reg342[(2'h3):(1'h1)]) >>> $signed(reg16))) >> ({($unsigned(wire356) >> {reg484,
                          reg491})} ?
                  (({reg475,
                      (8'hab)} != reg492[(3'h4):(1'h0)]) >>> reg483[(2'h2):(1'h0)]) : reg482[(2'h2):(2'h2)]));
              reg500 <= (($unsigned($unsigned((reg17 >= reg481))) ?
                  $signed(($signed(reg35) << forvar341)) : (($unsigned((8'hbf)) ^ (|reg457)) ?
                      $unsigned((&reg456)) : $unsigned($unsigned(reg497)))) > (reg352 >> $signed(reg468)));
            end
          else
            begin
              reg499 <= (reg22[(1'h0):(1'h0)] ^ ((((reg492 ?
                          reg321 : (8'hb5)) + forvar335[(1'h1):(1'h0)]) ?
                      (reg324[(4'h9):(2'h2)] > (reg492 | reg467)) : ($unsigned(forvar38) * (+(8'hbc)))) ?
                  $signed(($unsigned(reg345) ?
                      $unsigned(forvar474) : reg469[(1'h1):(1'h1)])) : (~|$signed((|reg42)))));
              reg500 = (reg36 ?
                  ((forvar485[(1'h0):(1'h0)] + $unsigned($signed(wire496))) ?
                      (((7'h43) ?
                          "DabS3zC9FT" : reg329) << {((7'h40) ~^ reg348)}) : {(-(reg332 ?
                              (8'hb9) : reg318))}) : ({$signed((wire453 <= forvar343))} ~^ {(!reg492),
                      (wire495 < $unsigned(reg497))}));
              reg501 = $unsigned({{$signed($unsigned(reg493)),
                      (&$signed(reg29))}});
            end
          for (forvar502 = (1'h0); (forvar502 < (1'h1)); forvar502 = (forvar502 + (1'h1)))
            begin
              reg503 <= (~&wire356);
              reg504 = (reg329[(3'h4):(2'h2)] ^ reg15[(3'h5):(2'h2)]);
              reg505 = (reg472 && reg34);
              reg506 <= ((~&wire9) & (reg332[(4'hb):(2'h3)] ^ $unsigned(reg477[(3'h4):(3'h4)])));
            end
          for (forvar507 = (1'h0); (forvar507 < (2'h2)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 = "lp7i99qUexzepU";
              reg509 = {$unsigned(((wire356[(3'h5):(1'h0)] ?
                          (~^forvar38) : reg345) ?
                      (8'ha3) : $signed((reg474 == reg486)))),
                  ((forvar507[(4'h8):(3'h5)] - reg338) >= $unsigned($signed((reg488 ?
                      reg466 : reg489))))};
            end
          reg510 <= (^~$signed($unsigned((~&$signed(reg462)))));
          if (((reg482 ? (^~$unsigned(reg482)) : forvar27) ?
              $unsigned((&(8'hae))) : reg338))
            begin
              reg511 = reg26;
              reg512 = reg331[(3'h7):(2'h3)];
              reg513 <= (8'hb1);
            end
          else
            begin
              reg511 = $unsigned((~|reg503[(4'hb):(1'h0)]));
            end
        end
      reg514 = reg463[(3'h7):(1'h0)];
    end
  assign wire515 = ((({$unsigned(reg34), (reg492 ? (8'ha0) : reg513)} ?
                           ((7'h42) ?
                               (+reg479) : (forvar315 << forvar22)) : (^~(&reg476))) ?
                       $signed((-reg486)) : ((~|$unsigned(reg505)) ?
                           ((reg506 >> reg462) ?
                               $unsigned(reg457) : (forvar470 ?
                                   reg36 : reg349)) : $unsigned((-reg503)))) | reg321[(2'h2):(1'h0)]);
  assign wire516 = reg461[(2'h2):(1'h0)];
  assign wire517 = {$unsigned($unsigned(((reg323 ? reg482 : (8'had)) ?
                           (reg482 == reg468) : (wire257 > reg24))))};
  always
    @(posedge clk) begin
      for (forvar518 = (1'h0); (forvar518 < (1'h1)); forvar518 = (forvar518 + (1'h1)))
        begin
          if ((reg512 * {((wire356[(4'hf):(4'hb)] ~^ {reg510}) ?
                  {(reg467 ? wire515 : wire517),
                      (reg316 ? reg28 : reg471)} : reg28[(1'h1):(1'h1)])}))
            begin
              reg519 <= reg41;
              reg520 <= ({reg458[(3'h5):(3'h4)],
                      $signed($signed((reg35 ? reg355 : (8'hac))))} ?
                  ((-(forvar317 && {reg482, forvar470})) ?
                      (reg33[(3'h4):(1'h0)] ?
                          (~|$signed(reg459)) : ((reg477 << reg508) ?
                              reg458[(2'h2):(1'h0)] : (reg462 > reg336))) : $unsigned((((8'hbf) ?
                              reg352 : reg332) ?
                          $unsigned(reg462) : (-forvar335)))) : $signed((8'ha9)));
            end
          else
            begin
              reg519 = (|{$unsigned(reg332[(1'h1):(1'h1)])});
            end
          for (forvar521 = (1'h0); (forvar521 < (3'h4)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 <= reg324[(5'h10):(2'h3)];
              reg523 <= reg16;
              reg524 <= {(~|(forvar351 ? {reg21} : $signed(reg17))),
                  "3XDlAKKVASsDT3zh5PN"};
            end
          reg525 <= $unsigned($signed({$signed(forvar470[(3'h5):(3'h4)]),
              (~|$unsigned(wire257))}));
          for (forvar526 = (1'h0); (forvar526 < (3'h4)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg527 = {($unsigned((reg474[(2'h3):(1'h1)] ~^ (^~wire357))) - {$signed("ScKzoBkb"),
                      "f2xaRWrYNJs"})};
              reg528 <= (forvar502[(2'h3):(2'h3)] <<< (($signed((~(8'hb7))) | ("PGm9dnW1YyaSvKIH1c" ?
                  wire517[(3'h4):(3'h4)] : (reg493 <<< reg465))) - forvar335));
            end
          for (forvar529 = (1'h0); (forvar529 < (1'h1)); forvar529 = (forvar529 + (1'h1)))
            begin
              reg530 <= (forvar459 >> $unsigned((((~reg474) ~^ $signed(reg24)) ^~ reg456[(2'h3):(1'h1)])));
              reg531 = $unsigned($signed(($unsigned($signed(forvar22)) ?
                  ({forvar20} <= reg348) : $signed((wire11 ?
                      reg345 : reg316)))));
            end
        end
      if ((!reg354[(2'h2):(1'h0)]))
        begin
          for (forvar532 = (1'h0); (forvar532 < (2'h3)); forvar532 = (forvar532 + (1'h1)))
            begin
              reg533 = $signed({"f6kfkhAqSO5"});
              reg534 <= (~|wire11[(2'h3):(1'h1)]);
            end
          for (forvar535 = (1'h0); (forvar535 < (1'h0)); forvar535 = (forvar535 + (1'h1)))
            begin
              reg536 <= wire496;
              reg537 <= (wire11[(4'hb):(3'h5)] ?
                  ((((~&reg487) ? reg31 : {(8'hbc)}) ?
                      (|(~|reg15)) : (&((8'ha0) * wire10))) - forvar526) : wire517);
              reg538 <= $signed({forvar521[(1'h0):(1'h0)]});
              reg539 = {wire257[(2'h2):(1'h0)]};
            end
          for (forvar540 = (1'h0); (forvar540 < (2'h2)); forvar540 = (forvar540 + (1'h1)))
            begin
              reg541 <= ($signed("dT1BVt") << reg33[(4'h8):(2'h2)]);
              reg542 = (reg338[(3'h4):(2'h3)] == forvar351);
              reg543 <= $unsigned(reg484);
              reg544 = ($signed(((|(reg472 ? wire515 : reg503)) ?
                      ((&reg13) > reg455) : ((|reg460) == $unsigned((8'hbf))))) ?
                  reg475 : ("4I5AI2" + {reg501}));
              reg545 <= "hZwk8SvZ6rgwp2";
            end
          reg546 <= {reg491,
              $signed({$signed($signed(wire257)),
                  (reg26 != "2CqJwfx7ldErIpiqbg")})};
        end
      else
        begin
          if (forvar532[(5'h10):(3'h6)])
            begin
              reg532 <= (-$unsigned(reg481));
              reg533 = ($signed(((|(reg527 < (8'ha1))) ?
                      (((8'ha8) <= reg494) ?
                          (reg348 == reg528) : forvar326) : ($unsigned(forvar314) ?
                          reg463 : (reg462 >>> reg42)))) ?
                  (({reg493[(3'h4):(2'h2)]} != reg347[(3'h7):(3'h7)]) - ((~&reg334[(4'h8):(2'h2)]) >>> $signed((reg25 && reg337)))) : reg355[(3'h6):(2'h3)]);
              reg534 <= $unsigned(($signed((!$unsigned(forvar502))) < (~^(+$signed(forvar326)))));
              reg535 <= ("KracwUk13zSiQHrf6hev" << wire312[(4'hb):(4'h8)]);
              reg536 = $signed(($unsigned((reg457 ?
                  {reg503} : $signed((8'ha4)))) > reg26[(4'hb):(4'ha)]));
            end
          else
            begin
              reg532 <= reg318;
              reg533 = $signed(forvar315[(1'h0):(1'h0)]);
              reg534 = {reg476[(3'h4):(1'h1)]};
            end
          if ((reg40[(1'h1):(1'h1)] ?
              ($signed(($signed(reg35) ^~ (^reg519))) ?
                  $signed(reg35) : {$signed((reg461 ? reg345 : (8'hb3))),
                      reg469}) : $unsigned($unsigned((~|$signed(wire312))))))
            begin
              reg537 <= (~|reg484[(1'h0):(1'h0)]);
              reg538 = $signed($unsigned((~|($unsigned(reg331) ?
                  (forvar343 >= (8'hbd)) : $signed(forvar351)))));
              reg539 = {$unsigned({(reg483 != {reg334})}),
                  {($unsigned({reg527, wire356}) ?
                          reg493 : (reg475 >= (|reg525)))}};
              reg540 <= $unsigned(($signed($unsigned(reg18)) ?
                  reg460[(3'h6):(2'h3)] : reg504));
              reg541 <= $unsigned($signed({$unsigned({(8'h9d), reg19}),
                  ($signed(forvar341) ^ forvar22[(4'h8):(3'h4)])}));
            end
          else
            begin
              reg537 <= reg505;
              reg538 = reg477[(2'h3):(1'h0)];
            end
          reg542 <= ($unsigned(($signed("iL9mUIhWZPgmyPGZhZ") ~^ (reg493[(3'h6):(2'h3)] ?
              (forvar518 != reg31) : forvar540))) >= $unsigned(reg533[(2'h2):(2'h2)]));
        end
      reg547 = ($signed($signed(reg349[(2'h3):(1'h1)])) ?
          ((forvar540 <<< $unsigned((reg532 ? reg461 : reg513))) ?
              (8'hb5) : (((reg324 >= reg500) ? {wire235} : forvar350) ?
                  reg456[(5'h10):(3'h4)] : {(reg478 ? wire495 : (8'hbd)),
                      $unsigned(forvar474)})) : ((~&(8'hac)) >> (reg467[(4'h9):(1'h1)] ?
              (~^(reg523 ? reg530 : reg34)) : $signed((reg21 ?
                  reg489 : reg538)))));
      reg548 <= reg337;
    end
  module358 modinst550 (.wire363(reg328), .wire360(forvar518), .wire359(reg514), .clk(clk), .y(wire549), .wire362(reg532), .wire361(reg494));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module358
#( parameter param451 = (({(|(^~(8'ha9))), ((!(8'hbc)) ? (8'hae) : ((8'hb0) ? (8'ha6) : (8'ha8)))} <<< ({{(8'ha4)}, (~&(8'hbb))} >>> (~^((8'hbc) ? (8'had) : (8'ha0))))) ? (|(~^(8'ha6))) : ((^(-((8'hba) | (8'hbe)))) ? (-(((8'had) ? (8'hbf) : (8'ha9)) == ((8'h9c) ? (7'h44) : (7'h42)))) : ((((8'hba) ^~ (8'ha5)) && (^~(8'hb7))) >= (~|(^~(8'hbe))))))
, parameter param452 = (^~({(8'h9e)} >>> (!param451))) )
(y, clk, wire363, wire362, wire361, wire360, wire359);
  output wire [(32'h436):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire363;
  input wire signed [(4'hf):(1'h0)] wire362;
  input wire signed [(4'hd):(1'h0)] wire361;
  input wire signed [(2'h3):(1'h0)] wire360;
  input wire signed [(5'h12):(1'h0)] wire359;
  reg signed [(4'hc):(1'h0)] reg450 = (1'h0);
  reg [(4'hd):(1'h0)] reg449 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg447 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar446 = (1'h0);
  reg [(4'hf):(1'h0)] reg445 = (1'h0);
  reg [(5'h12):(1'h0)] forvar444 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg443 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg441 = (1'h0);
  reg [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(4'ha):(1'h0)] reg439 = (1'h0);
  reg [(2'h2):(1'h0)] forvar438 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg435 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg434 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar432 = (1'h0);
  reg [(3'h6):(1'h0)] forvar431 = (1'h0);
  wire [(4'ha):(1'h0)] wire430;
  reg signed [(3'h5):(1'h0)] reg429 = (1'h0);
  reg [(4'h8):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg427 = (1'h0);
  reg [(3'h5):(1'h0)] forvar426 = (1'h0);
  reg [(4'ha):(1'h0)] forvar421 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar415 = (1'h0);
  reg [(4'ha):(1'h0)] reg425 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg424 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar423 = (1'h0);
  reg [(5'h15):(1'h0)] reg422 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg421 = (1'h0);
  reg [(3'h7):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg419 = (1'h0);
  reg [(4'hc):(1'h0)] reg418 = (1'h0);
  reg [(4'he):(1'h0)] reg417 = (1'h0);
  reg [(4'ha):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg415 = (1'h0);
  reg [(5'h13):(1'h0)] reg414 = (1'h0);
  reg [(4'hb):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar412 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg410 = (1'h0);
  reg [(4'h9):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar407 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg406 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg405 = (1'h0);
  reg [(5'h12):(1'h0)] forvar404 = (1'h0);
  reg [(5'h14):(1'h0)] forvar396 = (1'h0);
  reg [(5'h10):(1'h0)] forvar393 = (1'h0);
  reg [(3'h7):(1'h0)] reg392 = (1'h0);
  reg [(4'ha):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar402 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg401 = (1'h0);
  reg [(2'h2):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg398 = (1'h0);
  reg [(3'h7):(1'h0)] reg397 = (1'h0);
  reg [(5'h15):(1'h0)] reg396 = (1'h0);
  reg [(5'h14):(1'h0)] reg395 = (1'h0);
  reg [(2'h2):(1'h0)] reg394 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar392 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg391 = (1'h0);
  reg [(5'h12):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg389 = (1'h0);
  reg [(4'hb):(1'h0)] forvar388 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire387;
  reg [(4'he):(1'h0)] reg386 = (1'h0);
  reg [(4'h9):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg384 = (1'h0);
  reg [(4'ha):(1'h0)] reg383 = (1'h0);
  reg [(4'h9):(1'h0)] forvar382 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg381 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg380 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar379 = (1'h0);
  reg [(3'h5):(1'h0)] reg378 = (1'h0);
  reg [(5'h15):(1'h0)] reg377 = (1'h0);
  reg [(4'h9):(1'h0)] reg376 = (1'h0);
  reg [(5'h12):(1'h0)] reg375 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar374 = (1'h0);
  reg [(4'hb):(1'h0)] reg373 = (1'h0);
  reg [(4'ha):(1'h0)] forvar372 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg371 = (1'h0);
  reg [(3'h6):(1'h0)] reg370 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg369 = (1'h0);
  reg [(4'ha):(1'h0)] reg368 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg367 = (1'h0);
  reg [(5'h14):(1'h0)] forvar366 = (1'h0);
  reg [(2'h2):(1'h0)] forvar365 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg364 = (1'h0);
  assign y = {reg450,
                 reg449,
                 reg448,
                 reg447,
                 forvar446,
                 reg445,
                 forvar444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 forvar438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 forvar431,
                 wire430,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 forvar421,
                 forvar415,
                 reg425,
                 reg424,
                 forvar423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 forvar412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 reg405,
                 forvar404,
                 forvar396,
                 forvar393,
                 reg392,
                 reg403,
                 forvar402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 forvar392,
                 reg391,
                 reg390,
                 reg389,
                 forvar388,
                 wire387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 forvar379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 forvar374,
                 reg373,
                 forvar372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 forvar366,
                 forvar365,
                 reg364,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg364 = (^((~^wire361[(3'h6):(3'h4)]) ^~ wire361));
      for (forvar365 = (1'h0); (forvar365 < (3'h4)); forvar365 = (forvar365 + (1'h1)))
        begin
          for (forvar366 = (1'h0); (forvar366 < (1'h0)); forvar366 = (forvar366 + (1'h1)))
            begin
              reg367 = (wire361 ?
                  (!$unsigned((7'h42))) : wire361[(3'h5):(3'h5)]);
              reg368 <= wire362;
              reg369 <= wire359;
              reg370 = wire360;
              reg371 <= (-wire361);
            end
          for (forvar372 = (1'h0); (forvar372 < (3'h4)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 = ("" ?
                  {(~|({forvar366} ?
                          forvar372[(2'h3):(2'h3)] : reg370))} : $unsigned($signed($signed((~&forvar372)))));
            end
          for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
            begin
              reg375 <= forvar372[(4'ha):(2'h2)];
            end
          if ($signed({$signed($unsigned($signed(reg369)))}))
            begin
              reg376 = (($signed(reg373) | (forvar372[(3'h5):(1'h1)] ^~ forvar365[(1'h1):(1'h0)])) ?
                  (((^~forvar365) ?
                          (wire361[(4'h8):(2'h2)] >> {forvar372}) : ($unsigned(wire359) > (reg364 ?
                              wire359 : reg370))) ?
                      ((forvar366 >> (+reg373)) ?
                          reg367[(3'h6):(3'h5)] : reg375) : (-(-(-wire361)))) : forvar366[(3'h5):(3'h5)]);
              reg377 <= $unsigned(((~^reg368[(4'h9):(4'h9)]) ?
                  {(reg364[(4'h8):(3'h4)] ?
                          $signed((8'hab)) : (forvar366 ?
                              wire361 : (8'h9e)))} : reg367));
              reg378 <= $signed($unsigned($signed((^(&reg375)))));
            end
          else
            begin
              reg376 = $unsigned((&(~^(~|$signed(forvar365)))));
            end
          for (forvar379 = (1'h0); (forvar379 < (2'h3)); forvar379 = (forvar379 + (1'h1)))
            begin
              reg380 <= (~|wire360);
              reg381 <= reg370[(3'h4):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar382 = (1'h0); (forvar382 < (1'h1)); forvar382 = (forvar382 + (1'h1)))
        begin
          reg383 = ($unsigned("n2GFXE9z1KBtIY9DZJqv") << ((((wire360 ?
                  reg364 : reg377) * (wire360 ? reg375 : forvar374)) ?
              $signed(((8'hb1) ~^ forvar372)) : $unsigned($signed(forvar382))) ^~ {reg368,
              $unsigned({reg370, (7'h44)})}));
          reg384 = $unsigned((~|{$signed(forvar365[(1'h0):(1'h0)]),
              ((8'hbe) ~^ $unsigned(forvar365))}));
          reg385 <= $unsigned((8'haa));
        end
      reg386 = $signed($unsigned((8'ha0)));
    end
  assign wire387 = (~&$signed(((&(forvar379 ? reg383 : forvar366)) ?
                       wire359 : "ciGN06N1ECH")));
  always
    @(posedge clk) begin
      if ((+$unsigned((~&$signed((reg364 >> wire361))))))
        begin
          for (forvar388 = (1'h0); (forvar388 < (2'h2)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 <= {(!$unsigned(($signed(reg380) ?
                      (reg376 ? wire387 : wire360) : $signed(wire360))))};
              reg390 = ({($signed((reg384 ?
                      reg367 : forvar372)) ~^ $unsigned(reg384[(4'hd):(2'h3)]))} ^~ reg378[(2'h2):(1'h0)]);
            end
          reg391 <= $signed((forvar374 ?
              $unsigned((((8'hb7) ?
                  reg389 : forvar382) << $unsigned(forvar374))) : reg390));
          for (forvar392 = (1'h0); (forvar392 < (2'h2)); forvar392 = (forvar392 + (1'h1)))
            begin
              reg393 <= (-(!reg370));
              reg394 = $unsigned(reg364[(4'hb):(3'h5)]);
              reg395 <= (~^reg393[(3'h5):(1'h0)]);
              reg396 = ((~^(wire362[(4'hc):(2'h3)] ?
                  (reg377 ?
                      wire359 : $unsigned(reg391)) : wire359[(3'h5):(1'h1)])) > $unsigned(forvar365[(2'h2):(1'h1)]));
            end
          if (reg375[(5'h10):(1'h1)])
            begin
              reg397 = $signed((&"GSoCPRrz2whP"));
              reg398 <= (forvar365[(1'h1):(1'h0)] <<< reg369);
              reg399 <= ($signed($unsigned(({reg391, reg380} ?
                  (~|forvar392) : {wire362}))) != reg393[(3'h7):(2'h3)]);
              reg400 = (~"JUOt");
              reg401 <= (forvar366[(3'h5):(2'h2)] ?
                  $unsigned($signed(reg371[(4'h8):(2'h3)])) : $unsigned({((^~reg377) ?
                          (reg391 <<< (7'h43)) : {wire359})}));
            end
          else
            begin
              reg397 <= ($unsigned({$unsigned((8'hbe))}) ^ $unsigned($unsigned(("eHKq8u8RgsoPSPU9F" - ((7'h43) >> reg373)))));
            end
          for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
            begin
              reg403 = reg373[(3'h5):(1'h0)];
            end
        end
      else
        begin
          for (forvar388 = (1'h0); (forvar388 < (2'h3)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 = (^$unsigned((~&(~$signed(reg403)))));
              reg390 = reg395[(1'h0):(1'h0)];
              reg391 = $signed($signed((+(~(forvar392 < reg397)))));
            end
          reg392 = ($signed("iAvgDtB1Oac0ZECeeH") < reg373);
          for (forvar393 = (1'h0); (forvar393 < (3'h4)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 = (^{((~^((7'h43) ^~ forvar392)) ^~ wire362[(3'h4):(2'h3)]),
                  forvar374});
              reg395 <= (!{(!reg383)});
            end
          for (forvar396 = (1'h0); (forvar396 < (1'h0)); forvar396 = (forvar396 + (1'h1)))
            begin
              reg397 = reg399;
              reg398 = $unsigned((^$signed(reg383)));
            end
        end
      for (forvar404 = (1'h0); (forvar404 < (2'h3)); forvar404 = (forvar404 + (1'h1)))
        begin
          if (forvar382[(4'h8):(3'h5)])
            begin
              reg405 = $signed($unsigned($signed($unsigned({reg385}))));
              reg406 <= (^$unsigned({($unsigned(reg381) ?
                      (wire361 ? reg393 : wire360) : $unsigned(wire359)),
                  $unsigned($unsigned(forvar382))}));
            end
          else
            begin
              reg405 <= reg371;
            end
          for (forvar407 = (1'h0); (forvar407 < (3'h4)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 <= {$unsigned(reg401[(2'h2):(1'h0)])};
              reg409 <= {(~&{$signed(wire361[(1'h0):(1'h0)])}),
                  (-(($unsigned(forvar365) ?
                      (!reg376) : wire359) >= $unsigned($unsigned((8'ha6)))))};
              reg410 <= forvar404;
              reg411 <= reg391[(1'h1):(1'h1)];
            end
          for (forvar412 = (1'h0); (forvar412 < (2'h3)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 = forvar365[(1'h1):(1'h1)];
              reg414 <= $signed($unsigned($unsigned(($unsigned(reg395) & (forvar402 && reg370)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((~((reg391[(2'h2):(1'h1)] ?
          forvar393[(3'h4):(2'h3)] : $signed(reg397)) >= $signed((reg405 ^~ $unsigned(forvar407))))))
        begin
          if ((~&forvar379[(3'h6):(3'h5)]))
            begin
              reg415 <= $unsigned(forvar392);
              reg416 <= ($unsigned({{forvar379}, "g2DzM"}) ?
                  $signed((($unsigned(reg403) ?
                          (reg398 ? (8'ha0) : wire387) : (~^reg371)) ?
                      reg403[(3'h7):(3'h7)] : (reg386 & ((8'ha2) ?
                          reg377 : wire387)))) : $signed(wire360));
              reg417 = $signed("bpXPreY2YXi4CtNR");
              reg418 = reg384[(3'h5):(1'h0)];
            end
          else
            begin
              reg415 <= reg414;
              reg416 = (((8'ha0) || (^~reg364)) * $unsigned($unsigned({$unsigned(reg378)})));
            end
          if ((^~reg376))
            begin
              reg419 = forvar404[(1'h1):(1'h1)];
              reg420 = (reg403[(3'h6):(1'h0)] + forvar379);
              reg421 = reg380[(1'h0):(1'h0)];
            end
          else
            begin
              reg419 = {reg418};
              reg420 = (~|"MEa7L7KSB");
              reg421 = reg368;
              reg422 <= (reg394 ?
                  (wire363[(3'h6):(1'h1)] <<< $signed(reg400)) : $unsigned((7'h40)));
            end
          for (forvar423 = (1'h0); (forvar423 < (3'h4)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 <= $unsigned($signed({({(8'ha6),
                      reg408} <<< (reg392 ^~ (8'hb3))),
                  (~&$unsigned(reg406))}));
              reg425 <= $signed({reg369});
            end
        end
      else
        begin
          for (forvar415 = (1'h0); (forvar415 < (2'h3)); forvar415 = (forvar415 + (1'h1)))
            begin
              reg416 = (reg395 != {{(-wire360[(2'h2):(1'h0)]), forvar423}});
              reg417 <= (($unsigned((~&$unsigned((8'hae)))) ? reg367 : reg371) ?
                  (reg418[(1'h0):(1'h0)] ^ $signed((~^(~^reg398)))) : (+$signed($signed("I57qkGWozAtJdrZClzD"))));
              reg418 = $unsigned(forvar366[(5'h13):(5'h13)]);
              reg419 = {$signed(($signed($signed((8'hb2))) ?
                      ((+(8'hb8)) ?
                          reg377 : $signed(reg376)) : (-(reg411 && reg413)))),
                  reg419};
              reg420 <= reg389;
            end
          for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= ((-"YCKXFGaBP") != wire387[(2'h2):(1'h1)]);
            end
          for (forvar423 = (1'h0); (forvar423 < (1'h1)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 = ($signed($unsigned(reg421)) ? (~&(8'hb3)) : reg396);
              reg425 = ($signed(((8'hae) ?
                      $unsigned($signed((8'ha4))) : reg403[(4'h8):(3'h4)])) ?
                  ($signed(forvar396[(5'h13):(3'h4)]) ?
                      reg383[(4'h8):(3'h7)] : (-forvar365[(1'h0):(1'h0)])) : (+{(-(reg413 ?
                          forvar372 : wire361))}));
            end
          for (forvar426 = (1'h0); (forvar426 < (2'h2)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 = (~&forvar426[(3'h5):(2'h2)]);
              reg428 <= (+((~&((^reg376) + (forvar374 && reg410))) > (8'hbc)));
              reg429 = ($signed(forvar402) ?
                  (8'hae) : (reg400 <= (^(forvar379 >> reg408))));
            end
        end
    end
  assign wire430 = {(reg420 * ((reg427 ?
                               $unsigned(forvar402) : reg383[(3'h4):(1'h1)]) ?
                           reg401 : reg371))};
  always
    @(posedge clk) begin
      for (forvar431 = (1'h0); (forvar431 < (2'h3)); forvar431 = (forvar431 + (1'h1)))
        begin
          for (forvar432 = (1'h0); (forvar432 < (2'h2)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= reg420;
              reg434 = (~(reg408[(3'h4):(2'h2)] >>> forvar421[(4'h8):(1'h1)]));
              reg435 <= (~^reg381[(3'h7):(3'h7)]);
              reg436 <= ("mb00fO" ?
                  {$unsigned((reg386[(4'hd):(3'h6)] == ((8'hb4) * reg395))),
                      forvar431[(2'h2):(2'h2)]} : (~|reg417[(4'he):(4'h9)]));
            end
        end
    end
  always
    @(posedge clk) begin
      reg437 <= (forvar412 | $signed((reg420 ?
          "nDsHVtGwffXqCg0eXePz" : $signed(forvar365[(2'h2):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
        begin
          if ($signed((8'hb5)))
            begin
              reg439 = (((reg403 ?
                          ((reg410 ^ forvar388) * $signed(forvar402)) : {(!(8'hba))}) ?
                      $unsigned((^(~|(8'had)))) : (~&$signed((reg394 * forvar392)))) ?
                  $unsigned({reg427}) : $signed((8'ha5)));
              reg440 = (forvar382 && $unsigned($unsigned($signed((^~forvar426)))));
              reg441 = reg435;
            end
          else
            begin
              reg439 = ({{(forvar382 ?
                          reg418 : {(8'ha2)})}} >> $unsigned(({{reg401,
                          forvar382}} ?
                  reg410[(3'h4):(1'h0)] : (-{reg420}))));
              reg440 <= wire387;
              reg441 = (&"SMYdANGe8N6F0pao");
            end
          reg442 <= ((+"IItQ9TcQexYt") ? forvar407 : (8'hb1));
        end
    end
  always
    @(posedge clk) begin
      reg443 <= (((forvar404[(3'h6):(2'h3)] <<< forvar431) ?
          $signed(reg439[(4'h9):(2'h3)]) : reg396[(4'he):(4'ha)]) || reg413[(4'ha):(4'h8)]);
      for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
        begin
          reg445 <= reg394[(1'h0):(1'h0)];
          for (forvar446 = (1'h0); (forvar446 < (2'h2)); forvar446 = (forvar446 + (1'h1)))
            begin
              reg447 <= $signed(reg440[(1'h0):(1'h0)]);
              reg448 = (8'hbe);
            end
        end
      reg449 = forvar393[(3'h4):(2'h3)];
      reg450 <= (7'h43);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module259
#( parameter param310 = (((|((8'h9c) ? {(8'hb0), (8'hb5)} : ((8'hb8) ? (8'ha2) : (7'h40)))) ? (^~(((8'hb2) ^~ (8'hbe)) ? (+(8'hbf)) : ((8'h9e) ? (8'hbc) : (8'hb7)))) : (((~(8'hbb)) ? ((8'ha6) ? (8'ha1) : (7'h40)) : ((8'ha6) | (8'ha1))) - (~|{(8'h9c), (8'ha6)}))) ? (&{(((7'h41) >>> (8'hb8)) ? ((8'haa) ? (8'hbd) : (8'haf)) : {(8'hb3)})}) : (((^~{(8'h9e), (8'hb0)}) + (~|((8'h9d) - (8'ha9)))) - ((!(~^(8'hb3))) ? ({(8'hba)} | ((8'hb0) ? (8'ha0) : (8'hab))) : (8'h9f))))
, parameter param311 = {(param310 >= param310), param310} )
(y, clk, wire264, wire263, wire262, wire261, wire260);
  output wire [(32'h221):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire264;
  input wire [(4'ha):(1'h0)] wire263;
  input wire signed [(4'hc):(1'h0)] wire262;
  input wire [(3'h4):(1'h0)] wire261;
  input wire [(5'h15):(1'h0)] wire260;
  wire [(5'h14):(1'h0)] wire309;
  reg [(5'h10):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg307 = (1'h0);
  reg [(5'h10):(1'h0)] reg306 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg305 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg303 = (1'h0);
  reg [(3'h4):(1'h0)] forvar302 = (1'h0);
  reg [(5'h15):(1'h0)] reg301 = (1'h0);
  reg [(5'h11):(1'h0)] reg300 = (1'h0);
  reg [(3'h5):(1'h0)] reg299 = (1'h0);
  reg [(5'h13):(1'h0)] reg298 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar297 = (1'h0);
  reg [(4'he):(1'h0)] reg296 = (1'h0);
  reg [(3'h5):(1'h0)] reg295 = (1'h0);
  reg [(3'h4):(1'h0)] reg294 = (1'h0);
  reg [(4'h9):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar292 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg291 = (1'h0);
  reg [(3'h7):(1'h0)] reg290 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg287 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg286 = (1'h0);
  reg [(4'hf):(1'h0)] reg285 = (1'h0);
  reg [(4'hc):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar283 = (1'h0);
  reg [(4'hd):(1'h0)] reg282 = (1'h0);
  reg [(5'h12):(1'h0)] reg281 = (1'h0);
  reg [(5'h13):(1'h0)] forvar280 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar279 = (1'h0);
  wire [(3'h5):(1'h0)] wire278;
  reg [(4'hf):(1'h0)] reg277 = (1'h0);
  reg [(5'h13):(1'h0)] reg276 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg273 = (1'h0);
  reg [(5'h15):(1'h0)] forvar272 = (1'h0);
  reg [(4'he):(1'h0)] reg271 = (1'h0);
  reg [(5'h12):(1'h0)] reg270 = (1'h0);
  reg [(2'h2):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg267 = (1'h0);
  reg [(5'h15):(1'h0)] forvar266 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar265 = (1'h0);
  assign y = {wire309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 forvar302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 forvar292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 forvar280,
                 forvar279,
                 wire278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 forvar266,
                 forvar265,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar265 = (1'h0); (forvar265 < (1'h1)); forvar265 = (forvar265 + (1'h1)))
        begin
          for (forvar266 = (1'h0); (forvar266 < (1'h0)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 = wire260[(5'h13):(5'h13)];
              reg268 <= {(~^(~|(~^$unsigned(forvar265))))};
              reg269 = $signed(forvar266[(5'h15):(4'hb)]);
              reg270 <= (reg268 ?
                  {($signed("xr") * $signed((forvar265 ? forvar266 : (8'hb1)))),
                      (!((+(8'h9c)) + $unsigned(forvar265)))} : (^$signed(forvar265)));
              reg271 <= reg270[(5'h10):(1'h1)];
            end
          for (forvar272 = (1'h0); (forvar272 < (2'h2)); forvar272 = (forvar272 + (1'h1)))
            begin
              reg273 = ({(8'hb0),
                  $unsigned((wire263 >= reg267))} <= $signed($unsigned(reg268)));
              reg274 <= ((^$signed(wire264)) ?
                  $signed(reg269[(1'h0):(1'h0)]) : reg268);
            end
          if ($unsigned(forvar265))
            begin
              reg275 = (~&reg267);
            end
          else
            begin
              reg275 = wire264;
            end
          reg276 = forvar272;
          reg277 <= reg276[(4'hf):(4'ha)];
        end
    end
  assign wire278 = "J";
  always
    @(posedge clk) begin
      for (forvar279 = (1'h0); (forvar279 < (3'h4)); forvar279 = (forvar279 + (1'h1)))
        begin
          for (forvar280 = (1'h0); (forvar280 < (1'h1)); forvar280 = (forvar280 + (1'h1)))
            begin
              reg281 <= (forvar280 ?
                  reg267 : (-(forvar272 ?
                      $signed(wire260) : ({wire260} ~^ (&forvar280)))));
              reg282 = (reg275 ?
                  forvar272 : ({($unsigned((8'hb0)) + reg268)} | $signed(($unsigned((8'hb2)) ?
                      wire264 : forvar279))));
            end
          for (forvar283 = (1'h0); (forvar283 < (1'h1)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg284 = reg270;
              reg285 = reg274;
              reg286 <= $unsigned(((+(~^reg271)) < (forvar266[(2'h3):(2'h2)] != $signed((reg270 ?
                  forvar279 : reg284)))));
              reg287 <= $unsigned((((reg277[(4'h9):(3'h4)] - forvar266) ?
                      $signed(wire262) : forvar283) ?
                  (forvar280 <= reg284) : wire278));
            end
          reg288 = (($signed(reg285[(3'h4):(1'h0)]) << reg274[(3'h5):(2'h3)]) != ((~{$signed(forvar265),
              (wire264 ?
                  reg282 : reg270)}) && ((forvar279[(2'h2):(1'h0)] >= $unsigned(reg275)) ?
              ((forvar279 != forvar283) ?
                  $signed((8'hb4)) : (reg284 + reg287)) : (~$signed(forvar266)))));
          reg289 <= (!($unsigned({$unsigned((8'hae))}) ?
              reg288[(2'h3):(2'h2)] : "Ly46IU8M"));
          reg290 <= $signed($unsigned(wire261));
        end
      reg291 = reg269;
      for (forvar292 = (1'h0); (forvar292 < (1'h1)); forvar292 = (forvar292 + (1'h1)))
        begin
          if (reg284)
            begin
              reg293 = forvar272[(4'hd):(4'h8)];
              reg294 = reg275;
            end
          else
            begin
              reg293 <= forvar265;
              reg294 <= $unsigned({$unsigned((+reg281[(1'h1):(1'h0)]))});
              reg295 = (~reg274);
              reg296 = (|reg282);
            end
          for (forvar297 = (1'h0); (forvar297 < (1'h0)); forvar297 = (forvar297 + (1'h1)))
            begin
              reg298 = (((+$signed((+wire263))) ?
                  ($unsigned($unsigned(reg287)) <<< forvar272[(4'he):(4'h9)]) : $unsigned(forvar279[(1'h0):(1'h0)])) && "kSv92kKAY");
              reg299 <= wire262[(1'h0):(1'h0)];
            end
          reg300 = (^((8'h9f) < $unsigned(((+(8'hb2)) ^~ "xoNC9oekbkGs"))));
          reg301 = forvar283;
        end
      if ((({$signed("7gn1vUGC4YFWe6"),
                  ($unsigned(reg269) ? reg298 : (reg275 >> (8'hb4)))} ?
              (reg268 ~^ $signed($signed(forvar279))) : reg281) ?
          reg296 : ((^($signed(reg287) ?
              reg276[(5'h13):(4'h9)] : $unsigned(reg269))) ^~ (reg274[(2'h2):(1'h1)] ?
              ({reg298} ?
                  (wire262 || reg267) : $signed((8'ha3))) : $unsigned((reg284 ?
                  reg290 : reg301))))))
        begin
          for (forvar302 = (1'h0); (forvar302 < (2'h3)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg303 <= forvar283[(4'h9):(3'h4)];
              reg304 = forvar266;
              reg305 = $unsigned(reg290);
            end
        end
      else
        begin
          for (forvar302 = (1'h0); (forvar302 < (2'h2)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg303 <= wire263;
              reg304 <= forvar297[(3'h4):(1'h1)];
              reg305 <= $unsigned($unsigned((forvar292[(2'h3):(1'h0)] ?
                  (~^$unsigned(reg301)) : reg267[(4'h9):(3'h6)])));
              reg306 <= $unsigned($signed(forvar266[(5'h14):(4'h8)]));
            end
          reg307 <= {(+(((reg289 ?
                  reg306 : reg301) ~^ (|reg305)) != reg275[(1'h0):(1'h0)]))};
          reg308 <= reg294;
        end
    end
  assign wire309 = {{("BBVQx" >> forvar302[(2'h2):(1'h0)])}};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module239
#( parameter param256 = (~^{(&(((8'hbe) && (8'hb0)) ? (~|(8'hb2)) : {(8'hbb)})), (~(((8'hb4) - (7'h42)) <= ((7'h42) ? (8'ha6) : (8'hae))))}) )
(y, clk, wire243, wire242, wire241, wire240);
  output wire [(32'h7d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire243;
  input wire [(3'h4):(1'h0)] wire242;
  input wire [(4'hf):(1'h0)] wire241;
  input wire [(5'h10):(1'h0)] wire240;
  wire signed [(2'h2):(1'h0)] wire255;
  reg [(4'ha):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar253 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire252;
  reg [(4'ha):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg250 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg249 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar248 = (1'h0);
  wire [(3'h6):(1'h0)] wire247;
  wire signed [(5'h14):(1'h0)] wire246;
  wire [(3'h6):(1'h0)] wire245;
  wire [(4'hf):(1'h0)] wire244;
  assign y = {wire255,
                 reg254,
                 forvar253,
                 wire252,
                 reg251,
                 reg250,
                 reg249,
                 forvar248,
                 wire247,
                 wire246,
                 wire245,
                 wire244,
                 (1'h0)};
  assign wire244 = ((($signed((8'hbf)) ?
                       $unsigned((8'ha9)) : (wire243 <= "TKboJKJe")) <<< {{$signed(wire242)}}) <<< $signed(wire242[(1'h1):(1'h1)]));
  assign wire245 = (((((wire240 && wire240) ^ (wire240 >>> (7'h44))) ?
                               (+((8'ha6) ?
                                   wire240 : (8'ha4))) : wire242[(1'h1):(1'h1)]) ?
                           $signed("BCDlsfL8112k4") : (^~(+wire241))) ?
                       {(~(&$signed(wire241)))} : (~|(^wire240)));
  assign wire246 = ($signed($unsigned($signed(wire241))) == wire244);
  assign wire247 = (8'ha6);
  always
    @(posedge clk) begin
      for (forvar248 = (1'h0); (forvar248 < (2'h3)); forvar248 = (forvar248 + (1'h1)))
        begin
          reg249 = wire240[(5'h10):(2'h2)];
          if ((forvar248[(3'h7):(1'h1)] ? wire245 : "0EVHK87F98sWZ"))
            begin
              reg250 <= $unsigned(forvar248);
              reg251 = $signed((wire241[(3'h5):(1'h1)] && reg249[(1'h1):(1'h1)]));
            end
          else
            begin
              reg250 <= wire242;
              reg251 <= ((($signed(reg249[(1'h0):(1'h0)]) < (+(|wire247))) ?
                  {$signed(wire240),
                      $unsigned(wire243[(4'ha):(3'h6)])} : $unsigned((+$signed(forvar248)))) ~^ ($unsigned((^(reg251 << reg249))) & reg249[(2'h2):(1'h1)]));
            end
        end
    end
  assign wire252 = reg250;
  always
    @(posedge clk) begin
      for (forvar253 = (1'h0); (forvar253 < (3'h4)); forvar253 = (forvar253 + (1'h1)))
        begin
          reg254 = (reg250[(4'h8):(2'h3)] ?
              (wire241 ^ wire252) : ($unsigned(reg251[(1'h1):(1'h0)]) >= {forvar248,
                  ($signed(wire252) ? $unsigned((8'hba)) : "DTqZnDsG")}));
        end
    end
  assign wire255 = $unsigned($unsigned(forvar253));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module44
#( parameter param234 = (((!(~|(~(7'h42)))) ? (-(((8'hb3) || (8'ha1)) > ((8'h9e) > (8'hb3)))) : (((~&(8'hb7)) & (~(8'hb9))) ^~ (((8'hbb) ? (8'ha4) : (8'hbc)) ^ ((8'h9c) == (8'h9d))))) == (+(+(&(~(8'ha5)))))) )
(y, clk, wire49, wire48, wire47, wire46, wire45);
  output wire [(32'h832):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire49;
  input wire [(4'hc):(1'h0)] wire48;
  input wire signed [(5'h12):(1'h0)] wire47;
  input wire signed [(5'h11):(1'h0)] wire46;
  input wire signed [(3'h6):(1'h0)] wire45;
  wire [(5'h12):(1'h0)] wire233;
  reg [(2'h3):(1'h0)] reg232 = (1'h0);
  reg [(5'h10):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg230 = (1'h0);
  reg [(4'hc):(1'h0)] forvar229 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg228 = (1'h0);
  reg [(4'hc):(1'h0)] reg227 = (1'h0);
  reg [(5'h11):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg225 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg222 = (1'h0);
  reg [(5'h11):(1'h0)] reg221 = (1'h0);
  reg [(5'h11):(1'h0)] reg220 = (1'h0);
  reg [(4'he):(1'h0)] forvar219 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar218 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg216 = (1'h0);
  reg [(2'h3):(1'h0)] reg215 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg214 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg213 = (1'h0);
  reg signed [(4'he):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg211 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar210 = (1'h0);
  reg [(5'h15):(1'h0)] reg209 = (1'h0);
  reg [(5'h15):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg207 = (1'h0);
  reg [(3'h4):(1'h0)] reg206 = (1'h0);
  reg [(4'hb):(1'h0)] reg205 = (1'h0);
  reg signed [(4'he):(1'h0)] reg204 = (1'h0);
  reg [(2'h2):(1'h0)] reg203 = (1'h0);
  reg [(3'h6):(1'h0)] reg202 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg201 = (1'h0);
  reg [(3'h5):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg199 = (1'h0);
  reg [(5'h13):(1'h0)] forvar198 = (1'h0);
  reg [(4'hb):(1'h0)] forvar197 = (1'h0);
  reg [(3'h5):(1'h0)] reg196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg194 = (1'h0);
  reg [(3'h6):(1'h0)] reg193 = (1'h0);
  reg signed [(4'he):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar191 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg190 = (1'h0);
  reg [(3'h7):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg188 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg187 = (1'h0);
  reg [(5'h12):(1'h0)] reg186 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg185 = (1'h0);
  reg [(4'hc):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg183 = (1'h0);
  reg [(2'h2):(1'h0)] reg182 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg181 = (1'h0);
  reg [(5'h15):(1'h0)] reg180 = (1'h0);
  reg [(4'hf):(1'h0)] forvar179 = (1'h0);
  reg [(3'h7):(1'h0)] forvar178 = (1'h0);
  reg [(4'ha):(1'h0)] reg177 = (1'h0);
  reg [(4'he):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg175 = (1'h0);
  reg [(5'h12):(1'h0)] reg169 = (1'h0);
  reg [(5'h14):(1'h0)] forvar168 = (1'h0);
  reg [(5'h10):(1'h0)] forvar164 = (1'h0);
  reg [(5'h14):(1'h0)] reg174 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg173 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar169 = (1'h0);
  reg [(4'hb):(1'h0)] reg168 = (1'h0);
  reg [(4'h8):(1'h0)] reg167 = (1'h0);
  reg [(4'ha):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg163 = (1'h0);
  reg [(5'h10):(1'h0)] reg162 = (1'h0);
  reg [(5'h10):(1'h0)] forvar161 = (1'h0);
  reg [(3'h5):(1'h0)] reg160 = (1'h0);
  reg [(4'he):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar157 = (1'h0);
  reg [(5'h13):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg154 = (1'h0);
  reg [(4'ha):(1'h0)] forvar153 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg150 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg145 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar144 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire143;
  reg [(4'hb):(1'h0)] reg142 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar141 = (1'h0);
  reg [(3'h5):(1'h0)] reg140 = (1'h0);
  reg [(3'h7):(1'h0)] reg139 = (1'h0);
  reg [(4'he):(1'h0)] reg138 = (1'h0);
  reg [(4'hd):(1'h0)] reg137 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(5'h11):(1'h0)] forvar135 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar130 = (1'h0);
  reg [(4'hd):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg134 = (1'h0);
  reg [(5'h10):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg132 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg130 = (1'h0);
  reg [(5'h13):(1'h0)] reg129 = (1'h0);
  reg [(4'hb):(1'h0)] forvar128 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg127 = (1'h0);
  reg [(3'h5):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg125 = (1'h0);
  reg [(3'h4):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg123 = (1'h0);
  reg [(2'h2):(1'h0)] forvar122 = (1'h0);
  reg [(5'h15):(1'h0)] reg121 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg120 = (1'h0);
  reg [(5'h15):(1'h0)] reg119 = (1'h0);
  reg [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg117 = (1'h0);
  reg [(5'h13):(1'h0)] forvar116 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg114 = (1'h0);
  reg [(5'h11):(1'h0)] reg113 = (1'h0);
  reg [(3'h4):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg112 = (1'h0);
  reg [(4'hc):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg110 = (1'h0);
  reg [(5'h14):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar108 = (1'h0);
  reg [(5'h15):(1'h0)] reg107 = (1'h0);
  reg [(4'h8):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg105 = (1'h0);
  reg [(3'h7):(1'h0)] reg104 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar103 = (1'h0);
  reg [(5'h10):(1'h0)] reg102 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg100 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg99 = (1'h0);
  reg [(4'h8):(1'h0)] forvar98 = (1'h0);
  reg [(4'hf):(1'h0)] reg97 = (1'h0);
  reg [(4'hb):(1'h0)] reg96 = (1'h0);
  reg [(3'h7):(1'h0)] reg95 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg94 = (1'h0);
  reg [(3'h5):(1'h0)] forvar93 = (1'h0);
  reg [(4'hc):(1'h0)] reg92 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire91;
  wire signed [(4'h9):(1'h0)] wire90;
  reg [(2'h3):(1'h0)] reg89 = (1'h0);
  reg [(3'h6):(1'h0)] reg88 = (1'h0);
  reg [(5'h15):(1'h0)] forvar87 = (1'h0);
  reg [(2'h3):(1'h0)] forvar86 = (1'h0);
  reg [(4'he):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar84 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg83 = (1'h0);
  reg [(3'h7):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg81 = (1'h0);
  reg [(4'hc):(1'h0)] reg80 = (1'h0);
  reg [(4'he):(1'h0)] forvar79 = (1'h0);
  reg [(4'he):(1'h0)] forvar78 = (1'h0);
  reg [(5'h12):(1'h0)] reg77 = (1'h0);
  reg [(3'h6):(1'h0)] reg76 = (1'h0);
  reg [(4'hc):(1'h0)] reg75 = (1'h0);
  reg [(5'h12):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg73 = (1'h0);
  reg [(5'h13):(1'h0)] forvar72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg70 = (1'h0);
  reg signed [(4'he):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg68 = (1'h0);
  reg [(2'h2):(1'h0)] reg67 = (1'h0);
  reg [(3'h5):(1'h0)] forvar66 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg65 = (1'h0);
  reg [(5'h12):(1'h0)] reg64 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg62 = (1'h0);
  reg [(3'h4):(1'h0)] forvar61 = (1'h0);
  reg [(5'h13):(1'h0)] forvar60 = (1'h0);
  reg [(5'h15):(1'h0)] reg59 = (1'h0);
  reg [(4'hd):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg56 = (1'h0);
  reg [(3'h7):(1'h0)] forvar55 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg54 = (1'h0);
  reg [(5'h10):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg52 = (1'h0);
  reg [(2'h3):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar50 = (1'h0);
  assign y = {wire233,
                 reg232,
                 reg231,
                 reg230,
                 forvar229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 forvar218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 forvar198,
                 forvar197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 forvar179,
                 forvar178,
                 reg177,
                 reg176,
                 reg175,
                 reg169,
                 forvar168,
                 forvar164,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 forvar169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 forvar161,
                 reg160,
                 reg159,
                 reg158,
                 forvar157,
                 reg156,
                 reg155,
                 reg154,
                 forvar153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 forvar144,
                 wire143,
                 reg142,
                 forvar141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 forvar130,
                 reg128,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 forvar128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 forvar122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 forvar116,
                 forvar115,
                 reg114,
                 reg113,
                 reg108,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 forvar108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 forvar103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 forvar98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 forvar93,
                 reg92,
                 wire91,
                 wire90,
                 reg89,
                 reg88,
                 forvar87,
                 forvar86,
                 reg85,
                 forvar84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 forvar79,
                 forvar78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 forvar72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 forvar66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 forvar61,
                 forvar60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 forvar55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 forvar50,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar50 = (1'h0); (forvar50 < (2'h2)); forvar50 = (forvar50 + (1'h1)))
        begin
          if (forvar50)
            begin
              reg51 <= ((8'hac) ?
                  $signed((((wire48 ? (8'hb5) : wire47) ?
                      (forvar50 | (7'h43)) : $signed((8'ha1))) & ($unsigned((8'hbc)) ?
                      wire49[(4'h9):(4'h9)] : (wire48 ?
                          wire48 : wire47)))) : $unsigned($signed(wire47[(1'h0):(1'h0)])));
              reg52 <= ($signed((+wire49[(4'h9):(4'h9)])) ?
                  (~&(~&$signed((^wire45)))) : ($unsigned((forvar50 + ((8'hb3) > wire46))) || ({$signed(wire45),
                      wire45[(3'h6):(2'h2)]} * reg51[(2'h2):(1'h0)])));
              reg53 = (&wire47[(3'h7):(3'h4)]);
              reg54 = ((($unsigned((wire48 ? wire48 : reg52)) ?
                      wire48[(3'h6):(1'h1)] : (-(reg52 & reg53))) <= "d0Xlkp") ?
                  (+(({forvar50, reg52} ?
                      $unsigned(reg52) : $unsigned(wire48)) && (~wire45[(2'h3):(1'h0)]))) : $signed(((^$signed(wire45)) & ((forvar50 ?
                      forvar50 : reg53) >> $unsigned(reg52)))));
            end
          else
            begin
              reg51 <= $signed(($unsigned((^~wire46[(3'h4):(3'h4)])) || $unsigned($unsigned(wire49))));
              reg52 = reg53[(3'h6):(2'h2)];
            end
          for (forvar55 = (1'h0); (forvar55 < (1'h1)); forvar55 = (forvar55 + (1'h1)))
            begin
              reg56 <= $signed(wire49[(1'h0):(1'h0)]);
              reg57 = reg54[(2'h2):(2'h2)];
              reg58 <= wire46[(4'ha):(2'h2)];
              reg59 = reg58;
            end
        end
      for (forvar60 = (1'h0); (forvar60 < (2'h3)); forvar60 = (forvar60 + (1'h1)))
        begin
          for (forvar61 = (1'h0); (forvar61 < (1'h1)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 <= {(+$signed((reg57 ?
                      (reg51 + reg52) : (reg54 << reg53))))};
              reg63 = (($unsigned((7'h40)) >> reg51) ~^ reg59[(2'h3):(1'h1)]);
              reg64 = (forvar55[(3'h4):(3'h4)] ^ (((((8'hb1) << reg56) ?
                      (forvar50 == reg58) : reg59[(4'hc):(3'h7)]) != (+wire47)) ?
                  (~$signed((8'hbb))) : $unsigned($signed(forvar50[(2'h3):(2'h3)]))));
              reg65 <= (reg56 < (-((^~$signed(reg53)) ?
                  (8'ha6) : ($unsigned((8'ha8)) | $unsigned(wire49)))));
            end
          for (forvar66 = (1'h0); (forvar66 < (2'h3)); forvar66 = (forvar66 + (1'h1)))
            begin
              reg67 <= "Xm";
              reg68 = ($signed($signed((+(reg57 ?
                  reg51 : forvar55)))) < (|$signed({forvar60[(5'h12):(3'h4)]})));
              reg69 = (reg63 ?
                  wire48 : (reg53 ?
                      {reg59[(4'hf):(3'h7)]} : $signed(((reg58 >> forvar50) ?
                          forvar50 : $unsigned(reg53)))));
              reg70 = (+$unsigned(forvar66));
              reg71 = (("UMUdZJbZdko3t8bIBo1" <= (~^reg62[(3'h7):(3'h4)])) ?
                  ((forvar50 | (~|(^(8'hbb)))) == $unsigned($signed((^~(8'hb5))))) : ((($signed(forvar66) ?
                          $unsigned(forvar66) : (wire46 | reg59)) ?
                      reg62 : (reg69 >>> (~^reg65))) + $signed(("7nDDM" ?
                      wire47 : (reg68 ? (8'hab) : reg64)))));
            end
          for (forvar72 = (1'h0); (forvar72 < (3'h4)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 = (8'hb9);
              reg74 <= (8'hbc);
              reg75 = $unsigned((&$unsigned((+forvar61[(2'h3):(2'h2)]))));
              reg76 = ($unsigned((reg74[(4'h9):(1'h0)] < reg57[(1'h0):(1'h0)])) ?
                  ((~|(~$unsigned(reg71))) ?
                      $unsigned(((reg73 ? reg65 : (8'h9c)) ?
                          (forvar66 ?
                              (8'hb1) : forvar72) : ((8'hb0) - forvar55))) : $signed($signed($unsigned((8'ha7))))) : reg75[(3'h7):(3'h6)]);
            end
          reg77 = (&reg53[(3'h4):(2'h2)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar78 = (1'h0); (forvar78 < (1'h0)); forvar78 = (forvar78 + (1'h1)))
        begin
          for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 <= reg59;
              reg81 <= (8'hbd);
              reg82 = reg71[(3'h7):(2'h3)];
            end
          reg83 = $signed(reg59[(1'h0):(1'h0)]);
          for (forvar84 = (1'h0); (forvar84 < (1'h0)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 = $signed(((|reg57[(2'h3):(2'h2)]) > $unsigned($unsigned($unsigned(forvar50)))));
            end
        end
      for (forvar86 = (1'h0); (forvar86 < (1'h1)); forvar86 = (forvar86 + (1'h1)))
        begin
          for (forvar87 = (1'h0); (forvar87 < (1'h0)); forvar87 = (forvar87 + (1'h1)))
            begin
              reg88 = $signed(($unsigned((wire47[(5'h10):(4'hf)] == reg75[(4'h9):(3'h4)])) ?
                  forvar66 : $unsigned((reg76 ?
                      reg57 : (forvar84 ? reg85 : reg51)))));
            end
        end
      reg89 = ($signed(forvar50[(4'h8):(1'h1)]) - wire47);
    end
  assign wire90 = forvar61[(2'h3):(2'h3)];
  assign wire91 = $unsigned(((~$unsigned((reg51 ?
                      reg74 : wire49))) ^ forvar86));
  always
    @(posedge clk) begin
      reg92 <= reg64;
    end
  always
    @(posedge clk) begin
      for (forvar93 = (1'h0); (forvar93 < (2'h3)); forvar93 = (forvar93 + (1'h1)))
        begin
          if (forvar84)
            begin
              reg94 <= reg82[(3'h5):(3'h5)];
              reg95 <= {reg76[(3'h5):(3'h4)], wire47[(5'h11):(5'h11)]};
              reg96 = (((forvar50[(1'h0):(1'h0)] & $signed(forvar60[(4'hb):(3'h4)])) ?
                      $signed($unsigned(reg53[(3'h4):(3'h4)])) : (((~|reg64) ?
                          reg52 : (reg81 || reg58)) - $unsigned($signed(reg88)))) ?
                  (7'h43) : $unsigned((reg76 > $signed((reg77 >> (8'ha0))))));
            end
          else
            begin
              reg94 <= (|reg94);
              reg95 <= {reg85[(4'hc):(4'hc)]};
              reg96 = (8'h9c);
              reg97 = (+$signed((^~$signed(reg53[(4'ha):(4'h9)]))));
            end
          for (forvar98 = (1'h0); (forvar98 < (2'h3)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 = (reg65 <= {wire90,
                  $signed(((reg77 >>> wire47) < ((8'hb6) ? reg65 : reg58)))});
              reg100 = ({forvar55[(3'h5):(1'h0)]} ?
                  ($signed((8'hbc)) ?
                      reg65[(3'h4):(1'h1)] : {{(reg94 ~^ forvar61),
                              (reg99 << reg54)},
                          $unsigned({reg97})}) : (~^$unsigned({{forvar55,
                          reg59},
                      $signed(reg57)})));
              reg101 <= $unsigned((8'h9c));
            end
          reg102 <= (8'hb2);
        end
      if (reg53)
        begin
          for (forvar103 = (1'h0); (forvar103 < (2'h2)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 = ((8'hb6) << $signed((8'ha9)));
              reg105 = (8'hb0);
              reg106 = $signed($signed(reg82[(2'h3):(2'h2)]));
            end
          reg107 = reg76;
          for (forvar108 = (1'h0); (forvar108 < (3'h4)); forvar108 = (forvar108 + (1'h1)))
            begin
              reg109 <= $unsigned(($signed(reg106) ?
                  ($unsigned({reg81, reg104}) ?
                      $signed($signed(reg56)) : "D41CLDthQA") : (-$unsigned((~^wire47)))));
              reg110 <= $signed($unsigned($unsigned("qWrLpPx")));
              reg111 <= (((({(8'ha1),
                      forvar66} | reg100[(4'ha):(1'h0)]) && (~&(reg74 < reg89))) & ($unsigned((wire91 ?
                          reg94 : reg99)) ?
                      (8'hbd) : (~forvar55[(1'h1):(1'h0)]))) ?
                  {$signed((&wire48))} : $signed(reg59));
              reg112 = (reg80 <= $signed((^($signed(wire49) - reg77))));
            end
        end
      else
        begin
          for (forvar103 = (1'h0); (forvar103 < (1'h1)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 <= forvar66;
              reg105 <= $unsigned((reg92[(1'h0):(1'h0)] ?
                  $unsigned($unsigned((^reg75))) : ((8'hb0) ?
                      $unsigned((~|(8'hb5))) : (~^(reg105 ?
                          forvar72 : wire91)))));
            end
          if (((~&$signed($signed((reg56 > reg65)))) | reg71))
            begin
              reg106 <= (reg57[(1'h1):(1'h1)] ?
                  $unsigned((!({(8'ha3),
                      forvar60} | $unsigned(reg81)))) : ($unsigned({reg82[(2'h2):(1'h0)]}) ?
                      reg102[(3'h7):(3'h7)] : $signed(($signed(forvar72) - (reg110 ?
                          reg52 : (8'ha7))))));
              reg107 <= reg94[(1'h1):(1'h0)];
              reg108 = reg82[(3'h7):(2'h3)];
            end
          else
            begin
              reg106 <= ((reg58[(4'h9):(3'h4)] ~^ forvar84[(1'h1):(1'h0)]) ?
                  reg88 : ((~|{((8'hae) ^~ forvar87), reg106[(3'h4):(3'h4)]}) ?
                      reg71 : (8'had)));
              reg107 <= (reg80[(1'h1):(1'h1)] > {($unsigned($unsigned(reg94)) ?
                      (~|(forvar108 ? reg110 : reg109)) : $unsigned((8'h9f)))});
              reg108 <= (!(((^{reg105}) ?
                      (~(+(8'hae))) : reg59[(2'h3):(1'h1)]) ?
                  ({reg68[(3'h7):(2'h2)],
                      (|reg57)} ~^ reg52) : reg88[(2'h3):(2'h3)]));
            end
          if ($signed((forvar55 ?
              ($unsigned((reg69 || reg81)) ?
                  $signed((|reg54)) : reg101[(1'h1):(1'h1)]) : (~|({(8'ha3),
                      reg101} ?
                  (reg68 ^ (8'hba)) : $unsigned(wire45))))))
            begin
              reg109 = ((($signed($signed(wire90)) ?
                      ((reg107 ? reg54 : reg76) ?
                          (reg68 ?
                              reg70 : reg108) : $unsigned(reg65)) : ($signed(reg65) ?
                          (&forvar98) : forvar79)) & reg85) ?
                  (^(((8'h9c) * reg83) ?
                      $unsigned(forvar108) : (~"vY46AmiMcY"))) : $signed(forvar103));
              reg110 = wire90[(2'h2):(2'h2)];
              reg111 <= (~&reg106);
            end
          else
            begin
              reg109 <= $signed((($signed((reg88 && reg63)) ?
                      forvar78[(3'h6):(3'h4)] : reg108[(3'h4):(1'h1)]) ?
                  wire91 : $unsigned((forvar60[(4'he):(4'ha)] ?
                      $signed(reg56) : wire90))));
              reg110 <= ($signed(reg95) ?
                  reg96 : ($unsigned(reg82[(2'h2):(1'h1)]) ?
                      (^~(8'ha6)) : (^~{(reg105 ? reg88 : reg74)})));
              reg111 = reg51[(1'h1):(1'h1)];
              reg112 = ((^{reg80}) << $unsigned(reg97[(1'h1):(1'h1)]));
              reg113 = reg57[(1'h0):(1'h0)];
            end
          reg114 = {(!(((forvar86 ? forvar87 : reg65) == $signed((8'hac))) ?
                  (^~{(8'haa), reg106}) : (|$unsigned(reg95))))};
        end
      for (forvar115 = (1'h0); (forvar115 < (1'h0)); forvar115 = (forvar115 + (1'h1)))
        begin
          for (forvar116 = (1'h0); (forvar116 < (3'h4)); forvar116 = (forvar116 + (1'h1)))
            begin
              reg117 = $unsigned($unsigned($unsigned(reg95[(2'h3):(1'h0)])));
            end
          if (reg51[(1'h0):(1'h0)])
            begin
              reg118 <= reg107;
              reg119 = reg85;
              reg120 <= (-(~|forvar84));
            end
          else
            begin
              reg118 = reg117;
              reg119 = (reg53 >= ((~&(reg97[(4'h9):(3'h5)] <<< reg88)) >>> (+reg95[(2'h2):(1'h1)])));
              reg120 <= (8'ha6);
            end
        end
      reg121 = (-((~|wire48[(2'h2):(1'h1)]) >= reg120));
      for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
        begin
          reg123 <= $signed((+$unsigned((~|$unsigned((8'haf))))));
          reg124 = ($signed((reg107 ?
              ($unsigned(wire91) ?
                  (reg82 ~^ reg114) : $signed(wire46)) : ((~|reg63) ?
                  $signed((8'ha2)) : $signed(reg62)))) <<< ($signed(reg112[(2'h2):(1'h0)]) ?
              ((forvar86[(2'h2):(1'h0)] << (~wire91)) && (wire46[(1'h0):(1'h0)] ?
                  (wire49 ?
                      reg76 : wire47) : reg123)) : reg59[(5'h15):(5'h14)]));
          reg125 = (~({(wire46[(2'h3):(1'h0)] ? reg88 : (reg114 - (8'hb1)))} ?
              reg123 : $unsigned(forvar61)));
        end
    end
  always
    @(posedge clk) begin
      if (({reg106[(1'h1):(1'h1)]} - $unsigned((reg63[(3'h5):(2'h2)] == $signed($signed((8'h9d)))))))
        begin
          reg126 = wire49;
          reg127 <= $unsigned(reg69[(1'h0):(1'h0)]);
          for (forvar128 = (1'h0); (forvar128 < (1'h1)); forvar128 = (forvar128 + (1'h1)))
            begin
              reg129 <= ($signed($signed(reg81)) ?
                  reg113 : $signed(({(wire49 >= reg54)} ^ ((~|wire45) ?
                      reg106[(3'h4):(2'h2)] : reg123))));
            end
          reg130 = (~$signed(reg69[(2'h3):(1'h1)]));
          if ($signed($signed(reg59)))
            begin
              reg131 <= ($signed(reg85[(2'h3):(1'h0)]) >= reg121[(4'hf):(1'h0)]);
              reg132 = $unsigned($unsigned(((!reg124[(2'h2):(1'h1)]) ?
                  (8'ha1) : $unsigned((forvar72 ? reg59 : (8'ha2))))));
              reg133 = $signed({{"VZYAFmIrCSHI"}});
              reg134 <= reg107[(4'h8):(2'h2)];
            end
          else
            begin
              reg131 = (^~(($unsigned(wire49) ^~ "ubMBRK") ? reg124 : reg56));
              reg132 = (+forvar115[(1'h1):(1'h0)]);
              reg133 = (8'had);
              reg134 = reg70[(5'h10):(2'h3)];
            end
        end
      else
        begin
          reg126 = reg57[(1'h0):(1'h0)];
          if ((^~wire48[(1'h1):(1'h1)]))
            begin
              reg127 = (8'ha7);
              reg128 = $unsigned($unsigned((8'ha4)));
            end
          else
            begin
              reg127 = "tEGtpLWPaMCCM2";
              reg128 <= $signed((reg107 <<< $signed((wire47[(1'h1):(1'h0)] >> {reg95}))));
              reg129 <= (reg114 <<< "pcBbrPKESL84PbCszLoE");
            end
          for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= {(reg117 << (reg133 ?
                      forvar55 : (reg69[(2'h2):(2'h2)] ~^ (reg124 ?
                          reg133 : (8'haf)))))};
              reg132 = (~(^~"WbGZyHDuxmNaY7"));
              reg133 = $signed(reg106[(1'h0):(1'h0)]);
              reg134 <= ((~^(wire48 ?
                  reg114 : $signed((^~forvar84)))) || reg94);
            end
          for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= ((((8'haf) != (~$signed(forvar122))) ~^ (^~reg119[(1'h0):(1'h0)])) + $unsigned($signed($unsigned($unsigned(reg121)))));
              reg137 = reg111;
              reg138 = reg92[(4'hc):(3'h4)];
              reg139 <= (reg132 ?
                  reg75 : ((|(-(-forvar86))) ? (8'had) : (8'hbd)));
              reg140 = "0";
            end
          for (forvar141 = (1'h0); (forvar141 < (1'h1)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg142 = ($unsigned(($signed("WHFu25v") & $unsigned((&forvar135)))) ~^ (forvar78 ~^ ($unsigned($signed(reg108)) <= ((reg52 ?
                      forvar86 : reg54) ?
                  forvar60 : {reg83, reg125}))));
            end
        end
    end
  assign wire143 = $unsigned(($signed(wire47[(4'hb):(4'hb)]) ~^ (~&{(reg105 ?
                           reg108 : reg106)})));
  always
    @(posedge clk) begin
      if ({forvar141[(3'h6):(3'h4)]})
        begin
          for (forvar144 = (1'h0); (forvar144 < (1'h1)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 <= $signed($signed((-$signed($unsigned(reg111)))));
              reg146 = (^$unsigned($signed(($signed((8'hb7)) ?
                  ((8'hbf) >= reg107) : reg118))));
            end
          if ((!(~^(8'hae))))
            begin
              reg147 = ($signed($unsigned((~(&reg129)))) ^ reg101[(2'h2):(2'h2)]);
              reg148 <= $unsigned((!$signed(reg112)));
              reg149 = (~wire45[(2'h2):(1'h1)]);
              reg150 <= {(+wire90[(3'h5):(1'h1)])};
              reg151 = reg132[(1'h0):(1'h0)];
            end
          else
            begin
              reg147 = $signed("IU4G88r");
            end
          reg152 = {($unsigned(reg57) ?
                  reg130[(4'ha):(4'ha)] : (~^$unsigned($signed(forvar78))))};
          for (forvar153 = (1'h0); (forvar153 < (2'h3)); forvar153 = (forvar153 + (1'h1)))
            begin
              reg154 <= $signed(reg121[(5'h11):(4'he)]);
              reg155 <= reg77[(3'h7):(3'h4)];
              reg156 <= reg129[(4'hf):(4'h8)];
            end
        end
      else
        begin
          for (forvar144 = (1'h0); (forvar144 < (2'h2)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 = (8'hbc);
              reg146 = $signed(reg151[(3'h6):(3'h6)]);
              reg147 <= reg109[(1'h1):(1'h1)];
            end
        end
      for (forvar157 = (1'h0); (forvar157 < (1'h1)); forvar157 = (forvar157 + (1'h1)))
        begin
          reg158 = ((~|(reg51[(1'h0):(1'h0)] ?
                  $unsigned(forvar79) : ($signed(wire90) ? reg62 : reg101))) ?
              {reg123[(5'h10):(3'h7)],
                  (^reg96)} : $unsigned({{reg106[(2'h2):(1'h0)]},
                  reg138[(3'h6):(2'h2)]}));
          if ({((reg138 ? reg89 : reg137[(3'h6):(3'h4)]) ?
                  ((8'ha4) ?
                      forvar144 : (!$unsigned(reg63))) : forvar122[(2'h2):(1'h1)]),
              (reg146 & $signed(reg158[(4'ha):(3'h5)]))})
            begin
              reg159 = (reg134[(3'h6):(1'h0)] + (((!forvar135[(5'h11):(4'he)]) ^ ({(8'hae),
                      reg59} <= $signed(reg52))) ?
                  wire46 : (8'ha1)));
            end
          else
            begin
              reg159 <= $signed("r4nrk8IXes69Vy");
              reg160 = $signed((~|reg142));
            end
          for (forvar161 = (1'h0); (forvar161 < (2'h3)); forvar161 = (forvar161 + (1'h1)))
            begin
              reg162 <= (reg74 | ((($signed(reg75) ~^ "x") ?
                  ((reg131 && (7'h44)) == (^reg149)) : ($unsigned(wire45) < reg97[(4'hf):(1'h1)])) & $unsigned(reg154[(3'h5):(1'h1)])));
              reg163 = (~forvar98);
            end
        end
      if ($signed((reg51[(1'h0):(1'h0)] ?
          $unsigned(((~^forvar86) < $signed((8'hac)))) : $unsigned((!forvar157)))))
        begin
          if ($unsigned($signed(forvar84)))
            begin
              reg164 = $unsigned(((((reg57 ? (8'ha9) : reg105) ?
                  (reg105 || forvar93) : $unsigned(reg102)) && ($signed(reg155) ?
                  forvar122[(1'h1):(1'h1)] : $signed(forvar86))) & (!forvar72[(5'h11):(3'h5)])));
              reg165 = ((-reg96[(4'h9):(3'h6)]) * "Ona2D3fV4Hr");
              reg166 = reg162;
              reg167 = ($signed($unsigned(((reg148 >= reg139) ?
                  {reg53, reg147} : reg70))) & (^~reg112));
            end
          else
            begin
              reg164 = ((forvar66 & (-reg125)) ?
                  $signed({$unsigned({reg159, (7'h41)})}) : reg81);
              reg165 = ($unsigned((&((^~reg127) == {reg133}))) ^~ reg108[(2'h3):(1'h1)]);
            end
          reg168 <= $unsigned((+$unsigned(reg131)));
          for (forvar169 = (1'h0); (forvar169 < (2'h3)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg170 = $unsigned($unsigned(forvar128));
              reg171 <= {$signed(reg136), $unsigned(reg136[(2'h2):(1'h1)])};
              reg172 = (forvar50[(1'h0):(1'h0)] || reg80);
              reg173 = reg155;
            end
          reg174 = $signed(reg164);
        end
      else
        begin
          for (forvar164 = (1'h0); (forvar164 < (2'h2)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 = (~&forvar72);
              reg166 <= reg99;
            end
          reg167 = (-reg151);
          for (forvar168 = (1'h0); (forvar168 < (1'h0)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 <= ((((reg145 == $unsigned(reg160)) ?
                  forvar108[(5'h10):(4'hf)] : $unsigned((&reg74))) - ({reg158[(4'h8):(2'h2)]} ?
                  (~^wire143[(1'h1):(1'h0)]) : reg120)) + (forvar66 ^~ reg121));
              reg170 = {(~$unsigned($signed($unsigned(reg156))))};
            end
          if ({((reg82 ? $unsigned((8'haa)) : $signed($signed(reg164))) ?
                  reg112 : (+$signed(reg75[(2'h2):(1'h1)])))})
            begin
              reg171 <= (8'haa);
              reg172 <= (reg67 ? (&reg148) : reg57);
              reg173 = $signed({reg69, $signed(reg95[(2'h3):(2'h3)])});
              reg174 = reg139[(3'h6):(2'h2)];
              reg175 <= "nV0irmu";
            end
          else
            begin
              reg171 <= $unsigned(reg125);
              reg172 = $signed((8'hab));
              reg173 = $unsigned(reg67);
              reg174 <= reg149[(2'h2):(2'h2)];
            end
          reg176 = $unsigned(((($unsigned(reg69) ?
              wire48 : $signed(forvar87)) || "Js4951JsUwf") ^ $signed(reg108)));
        end
      reg177 = forvar116;
    end
  always
    @(posedge clk) begin
      for (forvar178 = (1'h0); (forvar178 < (1'h1)); forvar178 = (forvar178 + (1'h1)))
        begin
          for (forvar179 = (1'h0); (forvar179 < (2'h3)); forvar179 = (forvar179 + (1'h1)))
            begin
              reg180 <= (-$signed({reg131[(2'h3):(2'h2)]}));
              reg181 <= (~((~^(+(forvar108 ?
                  wire47 : (8'hbb)))) - $unsigned($signed((reg168 > reg69)))));
              reg182 = ($signed((8'had)) ?
                  ("" ?
                      forvar178 : (reg97 << (reg142[(4'h9):(3'h7)] | $signed(reg62)))) : $unsigned($signed($unsigned($signed(reg155)))));
              reg183 = (($signed(($unsigned(reg175) || $unsigned(reg129))) | reg96) < ((~^$unsigned($unsigned(reg145))) ?
                  reg129 : ((reg128[(2'h3):(1'h0)] - $signed(forvar179)) >> reg163[(3'h6):(3'h6)])));
            end
          reg184 = $unsigned(((!$signed(forvar55[(3'h7):(3'h7)])) > reg155[(3'h6):(1'h1)]));
          reg185 <= (($signed(($unsigned(reg65) ?
              $unsigned(reg177) : forvar141)) || {((forvar86 ?
                      reg102 : (8'hae)) ?
                  forvar122[(1'h0):(1'h0)] : reg131),
              (((8'hac) && reg53) ?
                  (forvar116 ?
                      reg174 : reg183) : $unsigned((8'ha7)))}) == "PLoQ2KVPe");
          if ($unsigned((!{({reg82} || reg131[(2'h3):(1'h1)])})))
            begin
              reg186 = reg53[(4'h8):(2'h3)];
              reg187 <= $signed((($signed((~|reg106)) & $signed((reg110 >> (8'ha5)))) ?
                  $signed(((forvar130 != forvar78) ?
                      (~reg74) : $signed(forvar157))) : {reg54, forvar168}));
              reg188 = forvar115;
              reg189 <= {(wire90 ? wire90 : (~|$unsigned($signed(reg152))))};
              reg190 = {($unsigned(reg111[(3'h5):(2'h3)]) ?
                      $signed($unsigned((!reg111))) : ($unsigned((forvar66 < forvar179)) < $signed(reg58[(4'ha):(2'h2)]))),
                  reg186};
            end
          else
            begin
              reg186 = $unsigned((^(^~$unsigned((+forvar179)))));
              reg187 <= (~reg139);
              reg188 = ($unsigned($unsigned("hfrftzE4aSPZ")) ?
                  forvar87[(3'h7):(3'h6)] : $signed($signed($unsigned(forvar168))));
              reg189 = $signed($signed(((-reg58) | $signed($signed((8'ha2))))));
              reg190 = (($unsigned(reg83[(1'h1):(1'h1)]) <<< ((!(reg156 <<< reg133)) ?
                      ((reg106 ?
                          wire46 : (8'haa)) <<< (|reg71)) : (forvar60[(5'h11):(1'h0)] ^~ reg123[(5'h12):(3'h6)]))) ?
                  $signed(($signed($unsigned(reg58)) ?
                      ((reg74 | (8'hb9)) > (reg169 <= reg127)) : {(reg168 ?
                              forvar60 : (8'ha6)),
                          {(8'hbd), reg133}})) : reg65);
            end
          for (forvar191 = (1'h0); (forvar191 < (1'h1)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 = $unsigned({($signed("aAe") >>> wire48[(4'ha):(4'h9)]),
                  {((8'ha9) <<< (reg174 != (8'ha0))),
                      ((wire90 ? forvar78 : reg100) << $signed(reg177))}});
              reg193 = $unsigned((^$unsigned(forvar153)));
              reg194 = (^~(~$signed((7'h43))));
              reg195 <= $signed(((($unsigned(reg95) + (forvar66 ^ reg76)) ?
                  (~&$signed(reg108)) : $signed((reg117 ?
                      reg123 : (8'hae)))) & $signed($signed($signed(reg151)))));
              reg196 = (($signed($signed(reg190[(3'h4):(2'h2)])) ?
                  "7zGXWXK" : ((reg180[(4'h9):(1'h1)] ?
                      $signed(reg131) : (reg148 ?
                          reg147 : reg68)) && (~(reg192 - reg100)))) >> reg52);
            end
        end
      for (forvar197 = (1'h0); (forvar197 < (2'h3)); forvar197 = (forvar197 + (1'h1)))
        begin
          for (forvar198 = (1'h0); (forvar198 < (2'h2)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= ({reg80[(4'h9):(3'h7)],
                      $signed($unsigned({reg187, forvar164}))} ?
                  $signed((+$signed({reg62}))) : reg83[(1'h1):(1'h0)]);
              reg200 <= $signed(reg173);
              reg201 = $unsigned({(~|"L9GMOZQbTh6DeUtmM5cl"),
                  {$signed((forvar66 ? reg193 : (8'ha7))), $unsigned(reg190)}});
              reg202 <= forvar144[(2'h3):(2'h2)];
              reg203 <= $signed($unsigned(((~reg167[(3'h7):(3'h6)]) < forvar108)));
            end
          reg204 = ($unsigned(forvar157) ?
              (~^reg156) : ((~&((reg168 ^ forvar128) & $unsigned(reg127))) && (!$unsigned((forvar164 ?
                  reg54 : wire47)))));
          reg205 <= (8'hb3);
          if ($signed($unsigned(((+(reg112 > reg201)) ?
              ((reg193 ? (8'h9d) : reg74) >> (~&forvar55)) : reg52))))
            begin
              reg206 <= forvar164[(4'hf):(3'h7)];
            end
          else
            begin
              reg206 = (!(~$signed(forvar103[(2'h3):(2'h2)])));
              reg207 = {(reg128[(4'hd):(2'h2)] ^ (({reg159} ?
                          (^~reg188) : forvar168) ?
                      (|$signed((8'had))) : $signed((forvar84 << wire49))))};
              reg208 <= $signed(($unsigned($unsigned(((8'hb0) ?
                      (8'hb9) : reg80))) ?
                  (reg136[(1'h0):(1'h0)] ?
                      forvar161[(2'h2):(1'h1)] : $signed($signed(reg162))) : forvar178[(1'h1):(1'h1)]));
              reg209 = ($unsigned((^~reg171[(4'hd):(4'hc)])) | $signed($signed((!((8'hab) && reg187)))));
            end
          for (forvar210 = (1'h0); (forvar210 < (1'h0)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= (^~reg150);
              reg212 = $signed((&(-{((8'ha2) << forvar103)})));
              reg213 <= reg200;
              reg214 <= reg129;
              reg215 = reg154;
            end
        end
      reg216 = $signed($signed(forvar55));
      reg217 = reg151;
      for (forvar218 = (1'h0); (forvar218 < (3'h4)); forvar218 = (forvar218 + (1'h1)))
        begin
          for (forvar219 = (1'h0); (forvar219 < (1'h0)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 <= $unsigned((~^reg119));
              reg221 <= {$signed($unsigned($unsigned((!forvar210)))),
                  $signed((reg139[(3'h5):(1'h0)] ?
                      ({(8'ha6)} || reg151[(1'h1):(1'h1)]) : ((reg181 ?
                          forvar116 : reg95) & reg155[(4'h9):(2'h2)])))};
              reg222 = (reg56 ? (+(8'ha2)) : reg163);
              reg223 = reg104;
              reg224 = {(((-reg140) <<< (^((8'hb0) ?
                      reg154 : reg172))) > $unsigned(((~|(8'hae)) ?
                      $unsigned(reg147) : ((8'hba) ? reg175 : reg64)))),
                  (forvar79 ? reg136 : reg175[(4'ha):(3'h6)])};
            end
          if (forvar197[(1'h1):(1'h1)])
            begin
              reg225 <= reg97[(3'h7):(1'h1)];
              reg226 = reg112;
              reg227 <= ((~&$unsigned((^(forvar164 == (8'h9f))))) != ($signed(reg200) ?
                  $unsigned(reg176[(4'hc):(4'ha)]) : $unsigned($unsigned(reg88))));
            end
          else
            begin
              reg225 = reg177;
              reg226 <= "C";
              reg227 = $unsigned((forvar218[(1'h0):(1'h0)] ^ (($signed(reg77) * ((8'hb1) ?
                  (8'hb5) : reg57)) | reg146)));
            end
          reg228 = $unsigned(forvar198[(1'h0):(1'h0)]);
          for (forvar229 = (1'h0); (forvar229 < (1'h1)); forvar229 = (forvar229 + (1'h1)))
            begin
              reg230 <= $signed((~&reg189));
              reg231 = $unsigned(($unsigned((^(reg70 ^~ (8'hbf)))) ?
                  (7'h42) : ($signed(reg81[(2'h3):(1'h1)]) ?
                      $signed((reg105 ?
                          (8'h9d) : wire48)) : (~$signed(reg112)))));
              reg232 <= {(+((reg224 ?
                      reg160[(2'h2):(2'h2)] : ((8'h9c) ?
                          reg64 : reg134)) >= (reg171[(4'ha):(3'h6)] & $unsigned(forvar103)))),
                  $signed(((|forvar178[(3'h5):(1'h0)]) ?
                      $unsigned(forvar122) : $signed($unsigned(wire46))))};
            end
        end
    end
  assign wire233 = $unsigned(((((reg105 & reg142) || $signed(reg67)) ?
                           $signed((8'hb4)) : (((8'hb9) ? reg126 : (8'hbf)) ?
                               $signed(reg180) : ((8'h9e) ?
                                   reg124 : forvar168))) ?
                       reg137 : reg63));
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h2f6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire3;
  input wire [(4'hc):(1'h0)] wire2;
  input wire signed [(2'h2):(1'h0)] wire1;
  input wire [(2'h3):(1'h0)] wire0;
  wire signed [(4'hd):(1'h0)] wire573;
  wire [(4'hc):(1'h0)] wire571;
  wire signed [(3'h6):(1'h0)] wire60;
  reg [(4'hb):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg58 = (1'h0);
  reg [(4'ha):(1'h0)] reg57 = (1'h0);
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg [(3'h6):(1'h0)] reg55 = (1'h0);
  reg [(2'h2):(1'h0)] reg54 = (1'h0);
  reg [(4'hc):(1'h0)] forvar53 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg52 = (1'h0);
  reg [(5'h11):(1'h0)] forvar51 = (1'h0);
  reg [(4'hf):(1'h0)] forvar50 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg48 = (1'h0);
  reg [(5'h15):(1'h0)] reg47 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg44 = (1'h0);
  reg [(4'h8):(1'h0)] forvar43 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar42 = (1'h0);
  wire [(4'h8):(1'h0)] wire41;
  wire [(5'h14):(1'h0)] wire40;
  reg signed [(5'h10):(1'h0)] reg39 = (1'h0);
  reg [(3'h6):(1'h0)] forvar29 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg37 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg34 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg32 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar31 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg26 = (1'h0);
  reg [(5'h10):(1'h0)] reg25 = (1'h0);
  reg [(5'h13):(1'h0)] forvar24 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg22 = (1'h0);
  reg [(4'hf):(1'h0)] reg21 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg20 = (1'h0);
  reg [(5'h12):(1'h0)] forvar19 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg17 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar12 = (1'h0);
  reg [(4'hf):(1'h0)] reg16 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg14 = (1'h0);
  reg [(4'h8):(1'h0)] reg13 = (1'h0);
  reg [(5'h15):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg11 = (1'h0);
  reg [(5'h12):(1'h0)] reg10 = (1'h0);
  reg [(2'h3):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg8 = (1'h0);
  reg [(4'hd):(1'h0)] reg7 = (1'h0);
  reg [(5'h12):(1'h0)] reg6 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4 = (1'h0);
  assign y = {wire573,
                 wire571,
                 wire60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 forvar53,
                 reg52,
                 forvar51,
                 forvar50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 forvar43,
                 forvar42,
                 wire41,
                 wire40,
                 reg39,
                 forvar29,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 forvar31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 forvar24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 forvar19,
                 reg18,
                 reg17,
                 forvar12,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 forvar5,
                 reg4,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 <= (~$signed(((+{wire1, wire0}) > (!wire3[(5'h14):(5'h13)]))));
      for (forvar5 = (1'h0); (forvar5 < (1'h1)); forvar5 = (forvar5 + (1'h1)))
        begin
          if ($unsigned(wire0))
            begin
              reg6 <= $signed("");
              reg7 = (^~$signed((8'hb4)));
            end
          else
            begin
              reg6 = {reg4[(2'h2):(1'h1)]};
            end
          if ((^(($signed($unsigned((8'hbf))) ?
              {wire3,
                  $signed(wire0)} : wire0[(2'h2):(2'h2)]) != "tgviOTXZPRLWi")))
            begin
              reg8 = ((($signed($signed(reg6)) ^ wire1) >= $signed(wire1[(2'h2):(2'h2)])) && wire3);
              reg9 = (&$signed(reg4));
            end
          else
            begin
              reg8 <= reg7[(4'ha):(2'h3)];
              reg9 = (&$signed($signed($unsigned(wire1[(1'h1):(1'h0)]))));
              reg10 <= wire1;
            end
        end
    end
  always
    @(posedge clk) begin
      reg11 = reg6;
      if ((+$unsigned({{reg11[(5'h10):(4'ha)]}})))
        begin
          reg12 = {(~^reg6), {(~forvar5)}};
          if ({forvar5})
            begin
              reg13 <= (^(reg11[(3'h4):(1'h1)] <<< (reg10 ?
                  reg11 : reg9[(2'h2):(1'h0)])));
              reg14 <= (reg12[(3'h4):(3'h4)] > $signed(($signed((-reg10)) ?
                  "n0sYKxoD7oF9XJ" : $unsigned($unsigned(reg11)))));
              reg15 = $signed({$signed(((reg6 <<< (8'ha5)) ?
                      $signed(reg11) : reg7[(2'h2):(1'h0)])),
                  ($signed({wire3}) - $signed((reg6 ? wire2 : wire2)))});
              reg16 = $unsigned($unsigned(reg15));
            end
          else
            begin
              reg13 = $unsigned(($unsigned($unsigned("Kg7fhJ")) ?
                  (^~"3JM4fVVJ3tkxIn") : reg14));
              reg14 = ($signed((({reg11} != (forvar5 >> reg9)) <<< wire1[(2'h2):(1'h0)])) ?
                  wire3 : $unsigned($signed(reg8)));
              reg15 <= (~|(~|(((|reg4) ?
                  {reg11, reg13} : (reg8 ?
                      (8'ha5) : wire2)) & reg15[(1'h1):(1'h1)])));
              reg16 <= ($signed(reg4) >>> reg4);
            end
        end
      else
        begin
          for (forvar12 = (1'h0); (forvar12 < (2'h2)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= ($signed($unsigned(reg13[(3'h7):(3'h6)])) ~^ $signed((|{"3PuNVPk2tN3Dq"})));
              reg14 <= {$signed(reg8[(4'he):(2'h3)]), reg4[(1'h1):(1'h0)]};
              reg15 <= wire1;
              reg16 = $unsigned(("ui4GKiJchyu18" < reg16));
              reg17 <= {({((wire2 > reg9) <<< $unsigned(reg4))} ?
                      forvar5 : {reg6, (8'hac)})};
            end
          reg18 <= (reg15 ? reg4[(4'h8):(1'h1)] : "735BJPu");
          for (forvar19 = (1'h0); (forvar19 < (2'h3)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 <= (!(^wire3[(5'h11):(3'h7)]));
              reg21 = (($signed((~$unsigned(reg4))) != (|($signed(reg15) ?
                      (~^(8'ha2)) : reg13[(2'h3):(2'h3)]))) ?
                  ((|$signed(reg8)) ?
                      reg16[(1'h1):(1'h0)] : $unsigned($signed({reg8}))) : (~&reg17[(2'h2):(2'h2)]));
              reg22 <= $unsigned($unsigned(reg7[(2'h3):(2'h3)]));
            end
        end
      reg23 <= {wire0[(1'h1):(1'h0)],
          {$unsigned(reg9),
              ($signed((^(8'hb8))) ?
                  (&((8'ha1) || (8'hb7))) : ((reg4 ? reg14 : reg4) ?
                      (8'hbc) : forvar19[(4'h9):(4'h9)]))}};
      if ($signed((($signed((reg11 ? reg18 : reg4)) ?
          reg23[(1'h0):(1'h0)] : $signed($signed(reg8))) && $signed({reg11[(1'h1):(1'h0)]}))))
        begin
          for (forvar24 = (1'h0); (forvar24 < (2'h2)); forvar24 = (forvar24 + (1'h1)))
            begin
              reg25 = (^~(((|{reg15, (8'h9f)}) ?
                      reg17 : (~|reg20[(3'h7):(3'h7)])) ?
                  $unsigned({reg17}) : (8'hb2)));
            end
          reg26 <= reg11;
          if ($signed(reg15))
            begin
              reg27 <= (reg12[(2'h2):(2'h2)] >>> (((~&{reg18}) ?
                  reg18[(3'h5):(2'h3)] : (|(^~reg16))) <<< reg4));
              reg28 <= $signed($unsigned({(^reg16), wire1}));
              reg29 = wire1[(1'h0):(1'h0)];
              reg30 = reg9;
            end
          else
            begin
              reg27 = (reg10[(3'h5):(2'h2)] ?
                  ((~reg9) >> $signed(({(8'h9d),
                      (8'hae)} == (|reg10)))) : forvar5[(1'h1):(1'h1)]);
              reg28 <= (|wire1);
              reg29 = ({$unsigned({(reg16 ? forvar19 : reg23)}),
                  wire2} <= reg4[(1'h1):(1'h0)]);
            end
          for (forvar31 = (1'h0); (forvar31 < (2'h3)); forvar31 = (forvar31 + (1'h1)))
            begin
              reg32 <= (($signed((~&$signed(reg30))) ?
                      {((reg28 ^ reg13) ?
                              (reg4 ?
                                  reg15 : reg27) : $unsigned(reg12))} : $unsigned(reg11[(4'hf):(1'h0)])) ?
                  $unsigned((reg23 > $signed(reg17[(1'h0):(1'h0)]))) : (^~(8'ha3)));
              reg33 <= ({(reg21 ?
                          (!(~&forvar5)) : $signed((wire0 ? reg15 : forvar5))),
                      reg8[(4'hf):(3'h6)]} ?
                  $signed(reg8) : $unsigned(forvar12));
              reg34 <= $signed(wire1);
            end
          if (reg33)
            begin
              reg35 = (~^$signed(forvar24[(4'hd):(4'ha)]));
              reg36 <= ((~&reg28) == (+((7'h43) || $signed($unsigned((8'ha9))))));
              reg37 = reg30;
              reg38 = $signed($unsigned($signed(reg29[(3'h5):(1'h1)])));
            end
          else
            begin
              reg35 = {{(((reg36 + reg6) ? {wire3} : (~^reg14)) ?
                          $signed(reg13) : (~|$signed(reg9)))},
                  $signed({$unsigned($signed(reg22))})};
              reg36 = reg16[(4'hc):(3'h5)];
              reg37 <= (~|(-forvar31));
              reg38 <= reg13;
            end
        end
      else
        begin
          for (forvar24 = (1'h0); (forvar24 < (1'h1)); forvar24 = (forvar24 + (1'h1)))
            begin
              reg25 <= forvar12[(1'h1):(1'h0)];
              reg26 <= reg22;
              reg27 = forvar5;
              reg28 <= $unsigned($unsigned({$unsigned(reg11)}));
            end
          for (forvar29 = (1'h0); (forvar29 < (1'h1)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 <= (((~($unsigned(reg22) ^~ reg14[(4'hd):(1'h1)])) ?
                  (reg29 ?
                      {$signed(reg27),
                          {reg29,
                              (8'ha7)}} : $unsigned(((8'ha5) ~^ reg25))) : ($signed((reg4 ?
                      reg16 : (8'hb9))) + (|(reg33 ?
                      reg38 : reg28)))) != reg29[(4'h8):(3'h5)]);
            end
        end
      reg39 <= (~&$unsigned(wire1));
    end
  assign wire40 = reg38;
  assign wire41 = {{reg38[(3'h6):(3'h5)]}};
  always
    @(posedge clk) begin
      for (forvar42 = (1'h0); (forvar42 < (2'h3)); forvar42 = (forvar42 + (1'h1)))
        begin
          for (forvar43 = (1'h0); (forvar43 < (3'h4)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg44 <= reg14;
              reg45 = ((!((forvar5[(2'h3):(1'h0)] ? $signed(reg8) : (~^reg12)) ?
                  ($signed(reg18) ?
                      $signed(reg25) : (reg38 > reg39)) : reg44)) ~^ (~|(8'hbb)));
              reg46 <= $unsigned($signed($unsigned(($signed(forvar42) ?
                  reg4 : wire2))));
            end
        end
      reg47 <= forvar19[(5'h12):(3'h4)];
      reg48 <= (((-$signed($signed(wire3))) ?
              $unsigned((~forvar43)) : (~^$unsigned(forvar19[(4'hd):(2'h3)]))) ?
          reg36[(3'h5):(2'h3)] : (reg26 ?
              $unsigned(reg30[(2'h2):(1'h0)]) : reg22));
      reg49 <= $signed($unsigned(reg23));
      for (forvar50 = (1'h0); (forvar50 < (2'h2)); forvar50 = (forvar50 + (1'h1)))
        begin
          for (forvar51 = (1'h0); (forvar51 < (1'h1)); forvar51 = (forvar51 + (1'h1)))
            begin
              reg52 <= $signed((^~($signed((~|reg13)) >>> {reg35})));
            end
          for (forvar53 = (1'h0); (forvar53 < (2'h3)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 = reg25[(2'h2):(2'h2)];
              reg55 <= $unsigned((8'haa));
              reg56 = reg45;
            end
          reg57 <= ($signed((((forvar43 ^~ (8'haa)) << (~&(7'h40))) >= (^$signed(forvar31)))) && $signed($unsigned($signed(((8'ha0) < reg4)))));
        end
    end
  always
    @(posedge clk) begin
      reg58 <= ($signed($unsigned((^~((8'hb7) >> reg25)))) >> {(~^$unsigned((forvar19 ?
              wire2 : reg49))),
          (+((forvar43 <<< (8'h9d)) ^~ forvar43[(3'h5):(2'h2)]))});
      reg59 <= forvar43[(3'h4):(1'h0)];
    end
  assign wire60 = ($signed((!(reg54[(1'h0):(1'h0)] ?
                      reg30 : (reg16 < wire40)))) << {{$unsigned(reg44[(3'h4):(2'h2)])},
                      (reg48 != $unsigned((wire0 ? (8'hb2) : reg4)))});
  module61 modinst572 (wire571, clk, forvar5, reg35, forvar50, reg34);
  assign wire573 = (^($signed(((reg25 * forvar19) <<< (-(8'had)))) ?
                       {reg45[(4'h9):(2'h2)]} : (reg34 * "o")));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module61  (y, clk, wire62, wire63, wire64, wire65);
  output wire [(32'h5c6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire62;
  input wire signed [(3'h7):(1'h0)] wire63;
  input wire [(4'h9):(1'h0)] wire64;
  input wire signed [(5'h15):(1'h0)] wire65;
  reg signed [(4'h8):(1'h0)] reg570 = (1'h0);
  reg [(4'h8):(1'h0)] reg569 = (1'h0);
  reg [(2'h2):(1'h0)] reg568 = (1'h0);
  reg [(4'h8):(1'h0)] reg567 = (1'h0);
  reg [(5'h15):(1'h0)] reg566 = (1'h0);
  reg [(4'hc):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar564 = (1'h0);
  reg [(5'h10):(1'h0)] reg563 = (1'h0);
  reg [(4'h8):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg561 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg560 = (1'h0);
  reg [(5'h10):(1'h0)] forvar559 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg558 = (1'h0);
  reg [(4'hf):(1'h0)] reg557 = (1'h0);
  reg [(2'h2):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg555 = (1'h0);
  reg [(5'h15):(1'h0)] forvar554 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg553 = (1'h0);
  reg [(4'hb):(1'h0)] forvar552 = (1'h0);
  wire signed [(4'he):(1'h0)] wire551;
  reg [(4'hb):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg548 = (1'h0);
  reg [(3'h5):(1'h0)] reg547 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar546 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg545 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar544 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg543 = (1'h0);
  reg [(2'h2):(1'h0)] reg542 = (1'h0);
  reg [(4'hc):(1'h0)] reg541 = (1'h0);
  reg [(4'hc):(1'h0)] forvar540 = (1'h0);
  reg [(3'h6):(1'h0)] reg539 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg538 = (1'h0);
  reg [(4'hf):(1'h0)] reg537 = (1'h0);
  reg [(5'h14):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg534 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar533 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar532 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg531 = (1'h0);
  reg [(3'h5):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg529 = (1'h0);
  reg [(2'h2):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg525 = (1'h0);
  reg [(3'h6):(1'h0)] forvar524 = (1'h0);
  reg [(5'h10):(1'h0)] reg523 = (1'h0);
  reg [(3'h6):(1'h0)] reg522 = (1'h0);
  reg [(5'h12):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar520 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg519 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg518 = (1'h0);
  reg [(3'h7):(1'h0)] reg517 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar516 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg515 = (1'h0);
  reg [(3'h7):(1'h0)] reg514 = (1'h0);
  reg [(2'h2):(1'h0)] reg513 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar512 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg511 = (1'h0);
  reg [(4'h9):(1'h0)] reg510 = (1'h0);
  reg [(3'h7):(1'h0)] reg509 = (1'h0);
  reg [(4'h9):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar507 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar506 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire476;
  wire [(4'hc):(1'h0)] wire263;
  wire signed [(4'hb):(1'h0)] wire66;
  reg signed [(5'h15):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg68 = (1'h0);
  reg [(5'h12):(1'h0)] reg69 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg71 = (1'h0);
  reg [(4'he):(1'h0)] reg72 = (1'h0);
  reg [(4'hb):(1'h0)] forvar67 = (1'h0);
  reg [(4'hf):(1'h0)] reg73 = (1'h0);
  reg [(2'h3):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg75 = (1'h0);
  reg [(3'h6):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg77 = (1'h0);
  wire [(3'h5):(1'h0)] wire78;
  wire signed [(5'h10):(1'h0)] wire79;
  wire [(3'h4):(1'h0)] wire80;
  reg signed [(3'h6):(1'h0)] forvar81 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg83 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar84 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg85 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg86 = (1'h0);
  reg [(3'h7):(1'h0)] reg87 = (1'h0);
  reg [(5'h14):(1'h0)] reg88 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg89 = (1'h0);
  reg [(3'h7):(1'h0)] reg90 = (1'h0);
  reg [(3'h6):(1'h0)] reg91 = (1'h0);
  reg [(5'h11):(1'h0)] reg92 = (1'h0);
  reg [(5'h15):(1'h0)] reg93 = (1'h0);
  reg [(4'hc):(1'h0)] reg94 = (1'h0);
  reg [(4'hb):(1'h0)] forvar95 = (1'h0);
  reg [(3'h7):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg98 = (1'h0);
  reg signed [(4'he):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg100 = (1'h0);
  reg [(5'h13):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar103 = (1'h0);
  reg [(4'h9):(1'h0)] reg104 = (1'h0);
  reg [(3'h5):(1'h0)] forvar89 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar92 = (1'h0);
  reg [(4'h9):(1'h0)] reg95 = (1'h0);
  wire [(4'h9):(1'h0)] wire105;
  wire signed [(2'h3):(1'h0)] wire106;
  wire [(4'hd):(1'h0)] wire107;
  wire [(4'hd):(1'h0)] wire108;
  wire [(5'h12):(1'h0)] wire109;
  reg [(2'h2):(1'h0)] forvar110 = (1'h0);
  reg [(3'h6):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg112 = (1'h0);
  reg [(4'hc):(1'h0)] forvar113 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar116 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg117 = (1'h0);
  reg [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg120 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg121 = (1'h0);
  reg [(4'hc):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar122 = (1'h0);
  reg [(4'ha):(1'h0)] reg123 = (1'h0);
  reg [(2'h3):(1'h0)] forvar124 = (1'h0);
  reg [(4'he):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg126 = (1'h0);
  reg [(3'h7):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg129 = (1'h0);
  reg [(3'h4):(1'h0)] reg130 = (1'h0);
  wire [(4'hb):(1'h0)] wire131;
  wire [(2'h2):(1'h0)] wire261;
  wire signed [(5'h12):(1'h0)] wire504;
  assign y = {reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 forvar564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 forvar559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 forvar554,
                 reg553,
                 forvar552,
                 wire551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 reg545,
                 forvar544,
                 reg543,
                 reg542,
                 reg541,
                 forvar540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 forvar533,
                 forvar532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 forvar524,
                 reg523,
                 reg522,
                 reg521,
                 forvar520,
                 reg519,
                 reg518,
                 reg517,
                 forvar516,
                 reg515,
                 reg514,
                 reg513,
                 forvar512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 forvar507,
                 forvar506,
                 wire476,
                 wire263,
                 wire66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 forvar67,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 wire78,
                 wire79,
                 wire80,
                 forvar81,
                 reg82,
                 reg83,
                 forvar84,
                 reg85,
                 reg86,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 reg94,
                 forvar95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 forvar103,
                 reg104,
                 forvar89,
                 forvar92,
                 reg95,
                 wire105,
                 wire106,
                 wire107,
                 wire108,
                 wire109,
                 forvar110,
                 reg111,
                 reg112,
                 forvar113,
                 reg114,
                 reg115,
                 forvar116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg110,
                 forvar122,
                 reg123,
                 forvar124,
                 reg125,
                 reg126,
                 reg127,
                 forvar128,
                 reg129,
                 reg130,
                 wire131,
                 wire261,
                 wire504,
                 (1'h0)};
  assign wire66 = (wire64 ^ {(!(+(|(8'ha9))))});
  always
    @(posedge clk) begin
      if (wire65[(4'he):(3'h4)])
        begin
          if (wire63[(1'h1):(1'h0)])
            begin
              reg67 <= (-($signed($unsigned((wire62 ? wire66 : wire65))) ?
                  $signed({wire66[(3'h4):(1'h0)]}) : (~|wire63)));
              reg68 = wire65;
              reg69 <= ($unsigned((~&$unsigned(wire66[(4'h9):(2'h2)]))) ?
                  wire64 : (((~|wire64[(3'h7):(3'h7)]) ?
                          $unsigned((wire62 <= reg67)) : wire62[(4'hc):(1'h1)]) ?
                      (^(wire63 ^ wire62[(2'h3):(2'h3)])) : (8'hb1)));
              reg70 = {((reg67 ?
                      ({wire66, (7'h43)} ?
                          (|wire65) : reg68) : wire66) != wire65)};
            end
          else
            begin
              reg67 <= (wire63[(3'h6):(2'h3)] ?
                  $signed(reg70) : ((+$unsigned(wire65)) >= (-(wire62 - reg68))));
              reg68 <= wire65[(4'ha):(1'h0)];
            end
          reg71 <= wire65;
          reg72 <= wire66;
        end
      else
        begin
          for (forvar67 = (1'h0); (forvar67 < (3'h4)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 = $unsigned($unsigned(($signed("hhh4vrsrG9GOLXCZ") - ((forvar67 ?
                      reg69 : wire62) ?
                  (reg69 ? reg71 : reg67) : reg67[(5'h15):(5'h15)]))));
              reg69 = reg72[(4'he):(4'he)];
              reg70 <= forvar67;
            end
          if ((^~{$signed($signed(wire64))}))
            begin
              reg71 <= (|reg68[(3'h7):(1'h1)]);
              reg72 = $unsigned((|(forvar67[(3'h6):(1'h0)] >>> reg69)));
              reg73 <= (~$signed(((reg69[(4'hb):(1'h1)] ?
                  reg70 : $signed(wire64)) != ((~|reg70) ?
                  ((8'ha8) ^ (8'ha9)) : $unsigned(reg69)))));
              reg74 = (reg73 * reg73[(1'h1):(1'h1)]);
            end
          else
            begin
              reg71 <= wire62;
              reg72 = reg71[(1'h0):(1'h0)];
              reg73 = $unsigned(($signed($unsigned((reg67 >> reg69))) ?
                  ($unsigned(reg67) ?
                      ($signed(reg68) > $unsigned((8'ha0))) : $signed((reg72 ?
                          reg74 : reg73))) : reg70[(3'h5):(1'h0)]));
              reg74 <= $signed((&($unsigned((reg74 ? (8'hb8) : reg72)) ?
                  (reg74[(1'h1):(1'h0)] ?
                      (&reg69) : reg69) : reg74[(1'h1):(1'h0)])));
              reg75 <= wire63[(1'h1):(1'h0)];
            end
        end
      reg76 = (-((|{$unsigned((8'h9e)), (-reg69)}) ?
          (((^~reg67) >= wire62[(4'hb):(2'h2)]) ?
              (|(reg72 ?
                  (7'h42) : forvar67)) : (~|$unsigned(forvar67))) : $signed({$signed(wire64)})));
      reg77 <= ((reg67[(4'he):(4'he)] ?
          {($unsigned(reg72) ~^ (!reg70))} : $signed($signed((reg76 ?
              reg69 : wire65)))) & (~&(($signed((8'hb9)) + (wire65 > (8'hab))) > $unsigned((~|reg73)))));
    end
  assign wire78 = ($unsigned((~|((reg76 ~^ wire65) >= ((8'ha8) && (8'hb6))))) != (8'hb9));
  assign wire79 = ((wire62[(2'h2):(1'h0)] <= $unsigned(reg70)) <= ({($signed(reg73) ?
                          (wire66 >>> reg77) : wire78)} <= reg77));
  assign wire80 = "s5XBR7N0GfDi8WraQg";
  always
    @(posedge clk) begin
      for (forvar81 = (1'h0); (forvar81 < (3'h4)); forvar81 = (forvar81 + (1'h1)))
        begin
          reg82 <= (8'ha2);
          reg83 <= (8'haa);
          for (forvar84 = (1'h0); (forvar84 < (1'h1)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 = ({reg73} * {$unsigned(($signed(wire62) ?
                      wire78[(3'h5):(1'h0)] : (&reg67))),
                  (^"dAb1e")});
              reg86 <= ((reg70[(3'h4):(1'h1)] ?
                  reg73 : reg85) <<< (~^"SidpD6LNZ8HVC8"));
              reg87 = ((^~wire63) ~^ "8t82HlaYipm");
              reg88 <= (($unsigned((((8'ha4) ? reg69 : reg68) ?
                      (reg85 ?
                          reg77 : (7'h44)) : (|wire64))) & (wire63 ^~ $signed(reg68[(4'hd):(1'h1)]))) ?
                  (reg87 ?
                      {(8'hb3),
                          reg69[(4'hb):(1'h0)]} : ((wire63[(3'h7):(3'h7)] | (|(8'hb3))) ?
                          wire79[(3'h6):(3'h5)] : ((&wire63) >> $signed((7'h44))))) : wire79);
            end
        end
      if ($signed(($signed(((~^reg76) ?
          reg68[(1'h1):(1'h1)] : wire79[(1'h0):(1'h0)])) == reg76[(3'h5):(1'h0)])))
        begin
          reg89 <= $unsigned($unsigned(((reg82[(1'h1):(1'h0)] ?
                  (reg88 ~^ reg75) : (reg67 ? forvar67 : wire80)) ?
              (~^(reg68 ~^ reg75)) : $unsigned($unsigned(reg72)))));
          if ((~^($signed($signed(forvar67[(3'h7):(2'h3)])) ?
              {{$signed(reg69)},
                  ($unsigned(reg67) >>> (reg73 ?
                      reg85 : (8'ha7)))} : {(^~((7'h44) ~^ reg73))})))
            begin
              reg90 <= {$signed(reg83)};
              reg91 <= wire65[(5'h10):(3'h5)];
              reg92 = reg89[(1'h1):(1'h1)];
              reg93 <= reg72;
              reg94 <= (&(|reg85[(2'h2):(2'h2)]));
            end
          else
            begin
              reg90 <= ((!(|reg91[(1'h0):(1'h0)])) ?
                  (&reg76) : ($unsigned(reg94[(3'h7):(3'h6)]) ?
                      $unsigned(((!(8'hac)) ?
                          reg94[(3'h6):(2'h3)] : $unsigned(reg82))) : $unsigned($signed(forvar84[(2'h2):(1'h1)]))));
              reg91 <= wire79;
              reg92 = (reg92 | (^$signed((-(reg85 ? reg68 : (8'hb3))))));
            end
          for (forvar95 = (1'h0); (forvar95 < (3'h4)); forvar95 = (forvar95 + (1'h1)))
            begin
              reg96 = ((+((|reg87[(3'h6):(3'h6)]) ?
                  reg91 : wire65[(5'h13):(3'h7)])) ^~ reg77[(4'h8):(4'h8)]);
              reg97 = {reg73[(4'h8):(2'h3)]};
            end
          if ($signed(reg90))
            begin
              reg98 = forvar95;
              reg99 <= (("hJ" ?
                  reg72[(4'h8):(3'h4)] : {$signed($unsigned(reg67)),
                      forvar67}) == $unsigned($unsigned($unsigned(reg82))));
              reg100 <= reg88[(4'hb):(3'h5)];
              reg101 = forvar84;
              reg102 = wire66[(2'h2):(1'h1)];
            end
          else
            begin
              reg98 = $signed(reg68);
            end
          for (forvar103 = (1'h0); (forvar103 < (2'h3)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 = (~^(((7'h42) ?
                  $unsigned($unsigned(reg98)) : (~^$signed(reg93))) && $signed($signed((reg77 * reg96)))));
            end
        end
      else
        begin
          for (forvar89 = (1'h0); (forvar89 < (2'h3)); forvar89 = (forvar89 + (1'h1)))
            begin
              reg90 <= $signed(reg82[(3'h6):(3'h6)]);
              reg91 = (wire78[(1'h1):(1'h0)] ?
                  (wire79 ^ (reg70[(2'h2):(2'h2)] ?
                      wire80 : (^(reg85 < wire65)))) : ($unsigned($signed((forvar103 * (7'h43)))) ?
                      (^~{reg98[(2'h2):(1'h0)]}) : ($unsigned((forvar84 ?
                              reg70 : reg88)) ?
                          $unsigned($unsigned(reg73)) : ($unsigned(wire65) < (+forvar81)))));
            end
          for (forvar92 = (1'h0); (forvar92 < (1'h0)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 = (8'h9e);
              reg94 = (reg70[(2'h3):(2'h2)] & $signed(($unsigned($unsigned((8'hba))) >= ((~|reg89) >> (wire65 ?
                  wire65 : reg87)))));
              reg95 <= {$unsigned(((~|(reg69 != reg97)) ?
                      $unsigned($signed(wire78)) : reg93))};
            end
        end
    end
  assign wire105 = reg100;
  assign wire106 = wire80;
  assign wire107 = ($signed(wire78[(3'h5):(1'h0)]) ?
                       reg97 : (($signed({reg82, forvar103}) ?
                               (~&reg77[(4'ha):(2'h2)]) : $signed(reg104)) ?
                           reg91[(2'h2):(1'h1)] : $unsigned($unsigned($unsigned((8'hb4))))));
  assign wire108 = (7'h44);
  assign wire109 = $signed((~&($unsigned(reg102[(4'hd):(4'hc)]) >>> reg77[(4'hf):(4'ha)])));
  always
    @(posedge clk) begin
      if (($unsigned($signed(((reg74 < reg68) ?
              $unsigned((7'h44)) : (reg68 ? reg85 : reg101)))) ?
          wire62 : {{($unsigned((7'h43)) ?
                      reg72[(4'hc):(3'h7)] : (reg99 ? (8'hb9) : reg91)),
                  $signed((wire107 ? reg83 : (7'h42)))}}))
        begin
          for (forvar110 = (1'h0); (forvar110 < (2'h3)); forvar110 = (forvar110 + (1'h1)))
            begin
              reg111 <= $signed((~&(^~"vz5h4Z0Q")));
              reg112 = (reg90 || ($signed(((~|reg101) || {wire64, wire64})) ?
                  ($signed(reg100) == reg104[(3'h5):(1'h1)]) : $signed({(&wire78)})));
            end
          for (forvar113 = (1'h0); (forvar113 < (1'h0)); forvar113 = (forvar113 + (1'h1)))
            begin
              reg114 = {(($unsigned((reg74 ? reg92 : wire63)) || ((reg76 ?
                              forvar92 : forvar110) ?
                          reg83[(1'h0):(1'h0)] : $signed(reg68))) ?
                      ((|$signed((8'ha4))) * wire64[(3'h7):(3'h4)]) : reg91),
                  $unsigned(reg71)};
              reg115 <= (((8'had) ?
                  (~$unsigned(((8'hbb) ?
                      forvar92 : reg114))) : reg90) < $unsigned(reg70[(4'h9):(1'h0)]));
            end
          for (forvar116 = (1'h0); (forvar116 < (2'h2)); forvar116 = (forvar116 + (1'h1)))
            begin
              reg117 <= forvar95;
              reg118 = $unsigned({(^~reg76), $signed({$unsigned(forvar81)})});
              reg119 = reg91[(3'h5):(2'h2)];
              reg120 = ((($signed((reg102 + reg89)) ?
                      ((7'h44) ?
                          (reg75 ?
                              wire62 : reg69) : $signed(reg83)) : $signed("RWLASRqecJl")) > reg67) ?
                  (^reg101[(4'h9):(2'h3)]) : ($signed($unsigned($signed(reg104))) ?
                      (^reg102) : ($signed((^forvar110)) ^~ forvar92[(1'h1):(1'h1)])));
            end
          reg121 = forvar92;
        end
      else
        begin
          reg110 = "bnQGp4CN";
        end
      for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
        begin
          reg123 <= (reg97[(4'ha):(3'h4)] ?
              $unsigned($unsigned((reg72 ? (+reg74) : reg110))) : reg68);
          for (forvar124 = (1'h0); (forvar124 < (2'h3)); forvar124 = (forvar124 + (1'h1)))
            begin
              reg125 <= (8'h9f);
              reg126 <= (~&$unsigned($unsigned((^~(reg121 ?
                  wire79 : reg100)))));
              reg127 <= {(~((~^reg67[(4'ha):(4'ha)]) ?
                      "E8v4k4z0sRXKWW" : ((~reg98) ?
                          wire79[(3'h4):(1'h1)] : reg115)))};
            end
          for (forvar128 = (1'h0); (forvar128 < (2'h3)); forvar128 = (forvar128 + (1'h1)))
            begin
              reg129 <= (&$signed(reg93));
            end
          reg130 = reg71;
        end
    end
  assign wire131 = $signed({(!($signed(reg77) >> (!reg90))),
                       (|$unsigned((+(8'hac))))});
  module132 modinst262 (wire261, clk, wire105, forvar92, forvar84, reg69, forvar128);
  assign wire263 = ($signed(((reg92[(2'h2):(1'h1)] ?
                               (8'hbc) : $signed(forvar103)) ?
                           (~&(reg110 ? wire108 : forvar95)) : ({wire66,
                                   reg94} ?
                               (reg130 ? reg99 : forvar116) : (forvar128 ?
                                   reg68 : (7'h43))))) ?
                       $signed(forvar110[(1'h1):(1'h1)]) : reg101);
  module264 modinst477 (.wire266(reg90), .wire265(reg73), .clk(clk), .wire267(reg120), .y(wire476), .wire269(reg77), .wire268(forvar103));
  module478 modinst505 (wire504, clk, wire108, reg93, reg82, wire131, reg72);
  always
    @(posedge clk) begin
      for (forvar506 = (1'h0); (forvar506 < (1'h1)); forvar506 = (forvar506 + (1'h1)))
        begin
          for (forvar507 = (1'h0); (forvar507 < (2'h3)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 <= forvar103[(4'ha):(2'h2)];
              reg509 <= (~^(^~$signed($signed(forvar506[(2'h2):(1'h0)]))));
              reg510 <= (((reg88 ?
                          forvar507[(4'hf):(1'h1)] : reg126[(3'h4):(1'h0)]) ?
                      reg98[(2'h3):(1'h1)] : forvar507[(5'h13):(3'h5)]) ?
                  $signed($unsigned("x7P")) : (!($signed($signed(reg126)) <= (^~$unsigned(wire65)))));
              reg511 = (reg73[(4'ha):(1'h1)] | wire106[(2'h3):(1'h0)]);
            end
          for (forvar512 = (1'h0); (forvar512 < (3'h4)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 <= $unsigned({(reg97[(1'h0):(1'h0)] != reg119),
                  $unsigned(reg95)});
              reg514 <= $signed({(~^$signed($signed(forvar122))),
                  ("YK0P" ?
                      {wire65[(5'h12):(4'h9)], (8'hbf)} : ({forvar122,
                          reg118} != $signed(wire476)))});
              reg515 <= ((&reg509) ~^ reg91);
            end
          for (forvar516 = (1'h0); (forvar516 < (2'h2)); forvar516 = (forvar516 + (1'h1)))
            begin
              reg517 <= forvar506;
              reg518 <= (!(((reg104 + reg87[(1'h1):(1'h1)]) << (wire106[(1'h1):(1'h0)] ^~ (~|reg71))) ?
                  reg74 : $unsigned((reg95[(3'h6):(1'h1)] ?
                      (reg129 << reg120) : reg82[(4'hb):(2'h3)]))));
              reg519 = {$signed($signed({reg92}))};
            end
          for (forvar520 = (1'h0); (forvar520 < (2'h3)); forvar520 = (forvar520 + (1'h1)))
            begin
              reg521 <= ($unsigned(((~&(reg515 ?
                  reg93 : (7'h40))) == (-$signed(forvar95)))) >= {(($unsigned(wire107) ?
                          $signed(wire261) : (&reg76)) ?
                      {reg111[(3'h4):(1'h1)]} : $signed((reg515 > (8'hbe))))});
              reg522 <= $signed((8'h9f));
              reg523 <= {reg110[(3'h5):(2'h2)], forvar122[(3'h6):(2'h3)]};
            end
        end
      for (forvar524 = (1'h0); (forvar524 < (1'h1)); forvar524 = (forvar524 + (1'h1)))
        begin
          reg525 <= (~&(reg75[(4'ha):(4'h8)] ?
              reg121[(2'h3):(2'h2)] : (&"sD6ms30FuQ")));
          if ((^~(reg519[(1'h0):(1'h0)] ?
              ($signed(wire131[(4'hb):(4'hb)]) ?
                  (~(reg121 >= (7'h42))) : $signed(reg67[(1'h1):(1'h0)])) : $unsigned(reg100[(2'h3):(2'h3)]))))
            begin
              reg526 <= reg71[(1'h0):(1'h0)];
              reg527 = ((8'hba) ^ reg74);
            end
          else
            begin
              reg526 <= {reg115};
              reg527 <= ((^~reg67[(3'h6):(2'h3)]) ?
                  {$unsigned(reg527),
                      (^reg117)} : $unsigned((("y" * {reg75}) > reg67[(5'h12):(3'h5)])));
              reg528 <= (+$unsigned($signed($unsigned(reg96[(3'h6):(1'h1)]))));
              reg529 = (|(forvar92[(3'h4):(1'h1)] != $unsigned({forvar95})));
            end
        end
      reg530 = ({$signed(forvar84)} < reg104);
      reg531 = $signed($unsigned(wire63));
      for (forvar532 = (1'h0); (forvar532 < (3'h4)); forvar532 = (forvar532 + (1'h1)))
        begin
          for (forvar533 = (1'h0); (forvar533 < (3'h4)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 <= {reg95[(3'h4):(2'h2)],
                  ({$unsigned((^~reg110)),
                      (^(forvar81 ? wire64 : reg118))} >= reg521)};
              reg535 <= $unsigned($unsigned($signed((|$unsigned(forvar103)))));
              reg536 <= $signed(((&(reg92 ^ {reg67})) ?
                  ($signed($unsigned((8'ha4))) ^~ (((8'hb7) <= forvar92) < ((8'hb6) ?
                      reg92 : (8'ha9)))) : reg111));
              reg537 <= $signed((&forvar89[(1'h0):(1'h0)]));
              reg538 = {$signed($unsigned(forvar89[(2'h3):(2'h2)])),
                  ($signed(((reg73 ? (8'ha4) : forvar516) ?
                      (reg125 | reg509) : (reg119 ?
                          reg86 : reg127))) < $signed(reg104))};
            end
          reg539 <= ($unsigned(reg70) ?
              ({($unsigned(reg518) ? (^reg99) : $signed(reg90))} ?
                  {reg83[(3'h7):(2'h2)],
                      wire62[(4'h8):(3'h6)]} : reg104) : {(~^((reg536 * forvar95) ~^ (~^wire107)))});
          for (forvar540 = (1'h0); (forvar540 < (1'h1)); forvar540 = (forvar540 + (1'h1)))
            begin
              reg541 <= $signed(reg82);
              reg542 <= ($unsigned(reg535) ?
                  $unsigned((reg95[(3'h4):(1'h1)] ^~ ((&wire64) ~^ (reg73 ?
                      (8'ha2) : (8'had))))) : (($unsigned((-reg508)) >>> (forvar84 & "9gcp6p")) ?
                      ({(reg541 <= wire63)} ^ (reg90 ?
                          (forvar124 != reg102) : (reg117 ?
                              forvar81 : reg71))) : $unsigned((8'ha1))));
              reg543 = (^(wire131 == {$signed($unsigned(reg526))}));
            end
          for (forvar544 = (1'h0); (forvar544 < (1'h0)); forvar544 = (forvar544 + (1'h1)))
            begin
              reg545 <= {reg508};
            end
          for (forvar546 = (1'h0); (forvar546 < (2'h3)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 <= $unsigned(reg89[(3'h5):(3'h4)]);
              reg548 = $unsigned($unsigned("KQ4qSnAxiIx"));
              reg549 <= $unsigned((&$unsigned($signed($unsigned(forvar512)))));
              reg550 <= wire64;
            end
        end
    end
  assign wire551 = (~reg91[(2'h3):(1'h0)]);
  always
    @(posedge clk) begin
      for (forvar552 = (1'h0); (forvar552 < (1'h0)); forvar552 = (forvar552 + (1'h1)))
        begin
          reg553 = (!(~^$signed(forvar128)));
          for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
            begin
              reg555 <= $signed((({{forvar544, (8'ha4)}} ?
                  $signed({reg86}) : (^~(reg542 && (8'hae)))) >= $unsigned($signed($unsigned(forvar124)))));
              reg556 <= $signed(($signed(forvar540[(4'hb):(1'h1)]) ?
                  ($signed({reg77, forvar533}) ?
                      ((reg88 << reg525) <<< $signed((7'h42))) : (&$signed(reg538))) : reg115));
              reg557 <= $unsigned($unsigned((^(wire504[(4'hc):(2'h3)] >= forvar516))));
              reg558 <= $unsigned((~&reg536[(4'he):(4'h9)]));
            end
          for (forvar559 = (1'h0); (forvar559 < (1'h0)); forvar559 = (forvar559 + (1'h1)))
            begin
              reg560 <= (^~({(wire109[(5'h10):(1'h1)] ? reg557 : (~|reg557))} ?
                  {"cz9te2IDzSib2gSW0MtV",
                      reg110[(2'h3):(1'h0)]} : reg531[(3'h4):(1'h0)]));
              reg561 <= reg94;
              reg562 = reg557;
              reg563 = reg92[(5'h10):(4'hc)];
            end
          for (forvar564 = (1'h0); (forvar564 < (2'h2)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 = {(wire504[(2'h3):(1'h1)] ?
                      forvar559[(4'hd):(3'h4)] : $unsigned(reg508))};
              reg566 <= (~^$unsigned((reg121[(1'h1):(1'h0)] ?
                  ((reg118 ? reg531 : reg96) ?
                      $signed(reg72) : forvar116[(3'h6):(3'h6)]) : $unsigned($unsigned((8'hb1))))));
              reg567 <= $unsigned(($unsigned("2JcPPGe5GJ") ?
                  "V8dfkm8T" : (($unsigned(reg86) ?
                          (~^reg90) : (reg537 ? reg75 : (8'ha6))) ?
                      $unsigned((reg555 ? (8'ha7) : reg543)) : (~|(reg543 ?
                          reg68 : reg114)))));
              reg568 <= reg100[(3'h5):(1'h0)];
              reg569 = reg531;
            end
        end
      reg570 = reg562[(2'h3):(1'h0)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module478
#( parameter param502 = ({(~&({(8'ha7), (8'ha8)} ^ ((8'hbe) ? (8'hbd) : (8'ha4)))), ((!{(8'hb5), (8'h9c)}) ? (((8'ha4) | (8'hbe)) == (7'h41)) : ((~^(7'h43)) ? ((8'ha8) >> (8'hb2)) : (+(8'hb3))))} ? (^~(((~|(8'hb9)) >= (&(8'ha3))) * ((-(8'hb7)) << (~^(8'hb0))))) : (-((((8'ha5) ? (7'h41) : (8'ha9)) ? (~&(8'hbc)) : {(8'hae)}) >> (~|{(8'hb5), (8'hbf)}))))
, parameter param503 = param502 )
(y, clk, wire483, wire482, wire481, wire480, wire479);
  output wire [(32'hc5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire483;
  input wire [(5'h13):(1'h0)] wire482;
  input wire signed [(5'h14):(1'h0)] wire481;
  input wire signed [(2'h2):(1'h0)] wire480;
  input wire signed [(4'h9):(1'h0)] wire479;
  wire [(5'h14):(1'h0)] wire501;
  wire signed [(4'hb):(1'h0)] wire500;
  wire [(5'h11):(1'h0)] wire499;
  wire signed [(2'h3):(1'h0)] wire498;
  wire signed [(2'h2):(1'h0)] wire497;
  reg signed [(5'h11):(1'h0)] reg496 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar494 = (1'h0);
  reg signed [(4'he):(1'h0)] reg493 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg491 = (1'h0);
  reg [(4'hc):(1'h0)] forvar490 = (1'h0);
  reg [(3'h5):(1'h0)] forvar489 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg488 = (1'h0);
  reg [(2'h2):(1'h0)] reg487 = (1'h0);
  reg [(5'h12):(1'h0)] forvar486 = (1'h0);
  reg [(2'h3):(1'h0)] reg485 = (1'h0);
  reg [(4'ha):(1'h0)] reg484 = (1'h0);
  assign y = {wire501,
                 wire500,
                 wire499,
                 wire498,
                 wire497,
                 reg496,
                 reg495,
                 forvar494,
                 reg493,
                 reg492,
                 reg491,
                 forvar490,
                 forvar489,
                 reg488,
                 reg487,
                 forvar486,
                 reg485,
                 reg484,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg484 <= $unsigned($unsigned(wire482));
      reg485 <= (wire481 ?
          wire483 : ($unsigned((~(wire481 ? wire482 : wire480))) ?
              (wire482 ?
                  (~^"offKwI") : (wire482[(4'h9):(4'h8)] ?
                      wire482 : $unsigned(wire479))) : (((wire482 ?
                      wire482 : (8'h9f)) ?
                  wire480[(1'h1):(1'h1)] : (wire482 ^~ (8'hbc))) <= (~^(wire482 < wire481)))));
      for (forvar486 = (1'h0); (forvar486 < (1'h0)); forvar486 = (forvar486 + (1'h1)))
        begin
          reg487 <= ($signed($signed($signed((wire482 <<< wire479)))) >= forvar486);
          reg488 = wire479;
        end
      for (forvar489 = (1'h0); (forvar489 < (2'h3)); forvar489 = (forvar489 + (1'h1)))
        begin
          for (forvar490 = (1'h0); (forvar490 < (2'h3)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 <= $signed((forvar490[(3'h7):(1'h0)] ?
                  $signed(($signed(forvar490) >>> reg484[(2'h3):(1'h0)])) : $signed("wSeBs9evk8SFou")));
              reg492 = ($unsigned($signed({wire483[(2'h2):(1'h1)],
                      (~&wire481)})) ?
                  $signed((|forvar490)) : (^$unsigned(wire483[(1'h0):(1'h0)])));
              reg493 <= (|reg488);
            end
          for (forvar494 = (1'h0); (forvar494 < (2'h3)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 = wire480[(2'h2):(2'h2)];
            end
        end
      reg496 = $unsigned({$signed($unsigned($signed(wire480))),
          forvar490[(4'ha):(2'h3)]});
    end
  assign wire497 = forvar494[(4'hd):(4'hb)];
  assign wire498 = wire483[(1'h1):(1'h1)];
  assign wire499 = (~($unsigned(wire498) ?
                       (forvar490 ?
                           $signed($unsigned(wire497)) : $signed("")) : $unsigned("G3kV0")));
  assign wire500 = wire481[(1'h1):(1'h1)];
  assign wire501 = wire482;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module264  (y, clk, wire269, wire268, wire267, wire266, wire265);
  output wire [(32'h9c9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire269;
  input wire signed [(4'hf):(1'h0)] wire268;
  input wire [(5'h10):(1'h0)] wire267;
  input wire [(3'h7):(1'h0)] wire266;
  input wire [(4'hf):(1'h0)] wire265;
  reg signed [(4'ha):(1'h0)] reg475 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg473 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg471 = (1'h0);
  reg [(3'h4):(1'h0)] reg470 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg469 = (1'h0);
  reg [(5'h15):(1'h0)] reg468 = (1'h0);
  reg [(4'hf):(1'h0)] reg467 = (1'h0);
  reg [(4'h8):(1'h0)] forvar466 = (1'h0);
  reg [(4'h8):(1'h0)] reg461 = (1'h0);
  reg [(3'h6):(1'h0)] reg465 = (1'h0);
  reg [(3'h4):(1'h0)] reg464 = (1'h0);
  reg [(4'hf):(1'h0)] reg463 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg462 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar461 = (1'h0);
  reg [(4'h8):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg459 = (1'h0);
  reg [(4'hc):(1'h0)] reg458 = (1'h0);
  reg [(5'h11):(1'h0)] reg457 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg456 = (1'h0);
  reg [(3'h5):(1'h0)] forvar455 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg453 = (1'h0);
  reg [(4'hc):(1'h0)] reg452 = (1'h0);
  reg [(5'h14):(1'h0)] forvar451 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg450 = (1'h0);
  reg [(4'h9):(1'h0)] forvar449 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg447 = (1'h0);
  reg [(5'h10):(1'h0)] reg446 = (1'h0);
  reg [(4'he):(1'h0)] reg445 = (1'h0);
  reg [(5'h15):(1'h0)] reg444 = (1'h0);
  reg [(5'h11):(1'h0)] forvar443 = (1'h0);
  reg [(5'h15):(1'h0)] reg442 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg440 = (1'h0);
  reg [(4'h9):(1'h0)] reg439 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg437 = (1'h0);
  reg [(2'h3):(1'h0)] reg436 = (1'h0);
  reg [(4'hb):(1'h0)] forvar435 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar433 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar432 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg430 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg429 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg428 = (1'h0);
  reg [(5'h10):(1'h0)] reg427 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar426 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg421 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg420 = (1'h0);
  reg [(4'hc):(1'h0)] forvar419 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg417 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar416 = (1'h0);
  reg [(5'h14):(1'h0)] reg415 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg412 = (1'h0);
  reg signed [(4'he):(1'h0)] reg411 = (1'h0);
  reg [(3'h5):(1'h0)] reg410 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar409 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar408 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg407 = (1'h0);
  reg [(3'h6):(1'h0)] reg406 = (1'h0);
  wire [(5'h14):(1'h0)] wire405;
  wire [(4'hf):(1'h0)] wire404;
  reg [(4'he):(1'h0)] reg403 = (1'h0);
  reg [(3'h5):(1'h0)] reg402 = (1'h0);
  reg [(3'h4):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg400 = (1'h0);
  reg [(3'h6):(1'h0)] reg399 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg398 = (1'h0);
  reg [(5'h11):(1'h0)] reg397 = (1'h0);
  reg [(2'h3):(1'h0)] forvar396 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg395 = (1'h0);
  reg [(3'h7):(1'h0)] reg394 = (1'h0);
  reg [(4'hd):(1'h0)] reg393 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar392 = (1'h0);
  reg [(5'h11):(1'h0)] reg391 = (1'h0);
  reg [(4'hf):(1'h0)] reg390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg387 = (1'h0);
  reg [(4'hb):(1'h0)] forvar386 = (1'h0);
  reg [(4'ha):(1'h0)] forvar385 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg383 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg382 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg380 = (1'h0);
  reg [(5'h12):(1'h0)] forvar379 = (1'h0);
  reg [(5'h12):(1'h0)] reg378 = (1'h0);
  reg [(3'h7):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg376 = (1'h0);
  reg [(3'h4):(1'h0)] forvar375 = (1'h0);
  reg [(4'he):(1'h0)] reg374 = (1'h0);
  reg [(3'h6):(1'h0)] reg373 = (1'h0);
  reg [(5'h12):(1'h0)] reg372 = (1'h0);
  reg [(3'h6):(1'h0)] reg371 = (1'h0);
  reg [(3'h5):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg369 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg368 = (1'h0);
  reg [(4'hb):(1'h0)] forvar367 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar366 = (1'h0);
  wire [(5'h14):(1'h0)] wire365;
  wire [(5'h11):(1'h0)] wire364;
  reg signed [(3'h4):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg361 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg360 = (1'h0);
  reg [(5'h12):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg358 = (1'h0);
  reg [(4'hb):(1'h0)] forvar357 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg356 = (1'h0);
  reg [(4'hd):(1'h0)] reg355 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg353 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar352 = (1'h0);
  reg [(3'h4):(1'h0)] forvar351 = (1'h0);
  reg [(3'h7):(1'h0)] reg350 = (1'h0);
  reg [(5'h15):(1'h0)] reg349 = (1'h0);
  reg [(3'h5):(1'h0)] reg348 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg347 = (1'h0);
  reg [(2'h2):(1'h0)] reg346 = (1'h0);
  reg [(2'h3):(1'h0)] forvar345 = (1'h0);
  reg [(4'hc):(1'h0)] reg344 = (1'h0);
  reg [(4'he):(1'h0)] reg343 = (1'h0);
  reg [(4'hc):(1'h0)] reg342 = (1'h0);
  reg [(4'h8):(1'h0)] forvar341 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar340 = (1'h0);
  wire [(5'h14):(1'h0)] wire339;
  reg [(5'h13):(1'h0)] reg338 = (1'h0);
  reg [(5'h12):(1'h0)] reg337 = (1'h0);
  reg [(4'ha):(1'h0)] reg336 = (1'h0);
  reg [(5'h13):(1'h0)] reg335 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg334 = (1'h0);
  reg [(5'h14):(1'h0)] reg333 = (1'h0);
  reg [(4'hc):(1'h0)] reg332 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar331 = (1'h0);
  reg [(5'h11):(1'h0)] forvar330 = (1'h0);
  reg [(5'h11):(1'h0)] reg329 = (1'h0);
  reg [(5'h11):(1'h0)] reg328 = (1'h0);
  wire [(4'h8):(1'h0)] wire327;
  reg [(4'h9):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar320 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg323 = (1'h0);
  reg [(3'h6):(1'h0)] reg322 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg320 = (1'h0);
  reg [(5'h11):(1'h0)] reg319 = (1'h0);
  reg [(3'h4):(1'h0)] reg318 = (1'h0);
  reg [(2'h2):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg316 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar315 = (1'h0);
  reg [(5'h14):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg313 = (1'h0);
  reg [(4'h9):(1'h0)] reg312 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg311 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg310 = (1'h0);
  reg [(4'h8):(1'h0)] reg309 = (1'h0);
  reg [(4'hb):(1'h0)] reg308 = (1'h0);
  reg [(4'hb):(1'h0)] reg307 = (1'h0);
  reg [(4'he):(1'h0)] reg306 = (1'h0);
  reg [(5'h14):(1'h0)] reg305 = (1'h0);
  reg [(2'h3):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg303 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg299 = (1'h0);
  reg [(5'h10):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar297 = (1'h0);
  reg signed [(4'he):(1'h0)] reg296 = (1'h0);
  reg [(4'hf):(1'h0)] reg295 = (1'h0);
  reg [(3'h5):(1'h0)] reg294 = (1'h0);
  reg [(5'h13):(1'h0)] reg293 = (1'h0);
  reg [(2'h2):(1'h0)] reg292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg291 = (1'h0);
  reg [(4'he):(1'h0)] forvar290 = (1'h0);
  reg [(2'h3):(1'h0)] reg289 = (1'h0);
  reg [(5'h14):(1'h0)] reg288 = (1'h0);
  reg [(5'h15):(1'h0)] reg287 = (1'h0);
  reg [(5'h11):(1'h0)] reg286 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg284 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar283 = (1'h0);
  reg [(4'h8):(1'h0)] reg282 = (1'h0);
  reg [(5'h15):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg280 = (1'h0);
  reg [(4'hb):(1'h0)] reg279 = (1'h0);
  reg [(5'h11):(1'h0)] forvar278 = (1'h0);
  reg [(4'hd):(1'h0)] reg277 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar276 = (1'h0);
  reg [(5'h15):(1'h0)] reg275 = (1'h0);
  reg [(4'he):(1'h0)] reg274 = (1'h0);
  reg [(3'h7):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg272 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar271 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire270;
  assign y = {reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 forvar466,
                 reg461,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 forvar461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 forvar455,
                 reg454,
                 reg453,
                 reg452,
                 forvar451,
                 reg450,
                 forvar449,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 forvar443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 forvar435,
                 reg434,
                 forvar433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 forvar419,
                 reg418,
                 reg417,
                 forvar416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 forvar409,
                 forvar408,
                 reg407,
                 reg406,
                 wire405,
                 wire404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 forvar396,
                 reg395,
                 reg394,
                 reg393,
                 forvar392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 forvar386,
                 forvar385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 forvar379,
                 reg378,
                 reg377,
                 reg376,
                 forvar375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 forvar367,
                 forvar366,
                 wire365,
                 wire364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 forvar357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 forvar352,
                 forvar351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 forvar345,
                 reg344,
                 reg343,
                 reg342,
                 forvar341,
                 forvar340,
                 wire339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 forvar331,
                 forvar330,
                 reg329,
                 reg328,
                 wire327,
                 reg326,
                 forvar320,
                 forvar317,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 forvar315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 forvar290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 forvar278,
                 reg277,
                 forvar276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 forvar271,
                 wire270,
                 (1'h0)};
  assign wire270 = $unsigned(($signed((wire268 ^ wire266[(2'h3):(1'h1)])) >> ((~^wire266) - $unsigned((^(8'hb9))))));
  always
    @(posedge clk) begin
      for (forvar271 = (1'h0); (forvar271 < (3'h4)); forvar271 = (forvar271 + (1'h1)))
        begin
          if ((wire268 - $unsigned(wire266)))
            begin
              reg272 = $unsigned((((~|(~&wire265)) ?
                  $unsigned((wire269 ?
                      forvar271 : wire270)) : $unsigned((wire265 ?
                      wire270 : wire268))) - forvar271));
            end
          else
            begin
              reg272 <= {((wire268 ?
                          $unsigned((forvar271 ^~ wire268)) : (!$signed(wire266))) ?
                      $unsigned((+$signed((8'hb6)))) : "U6")};
              reg273 = wire265[(1'h1):(1'h0)];
              reg274 = wire267;
            end
        end
      reg275 <= {forvar271, wire270[(1'h0):(1'h0)]};
      for (forvar276 = (1'h0); (forvar276 < (1'h0)); forvar276 = (forvar276 + (1'h1)))
        begin
          reg277 = $unsigned((8'ha9));
          for (forvar278 = (1'h0); (forvar278 < (1'h0)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= $unsigned($signed({"W4"}));
              reg280 <= {(+(((~^wire265) > reg279) >>> (|$unsigned(forvar278)))),
                  $unsigned($signed(wire268[(3'h7):(2'h2)]))};
              reg281 <= reg277[(3'h7):(2'h2)];
              reg282 <= ($signed($unsigned((~{reg277}))) ?
                  (reg277[(3'h6):(2'h3)] ?
                      reg272 : $signed(wire269[(1'h0):(1'h0)])) : (reg272[(3'h6):(3'h4)] ?
                      ($signed((wire265 | (8'ha7))) ?
                          $unsigned((wire268 > wire267)) : $unsigned((~^reg277))) : forvar278[(4'hc):(4'hb)]));
            end
        end
      for (forvar283 = (1'h0); (forvar283 < (3'h4)); forvar283 = (forvar283 + (1'h1)))
        begin
          reg284 <= reg274;
          if ((($signed((~&"SNK5")) ~^ ($unsigned((wire270 ?
              reg274 : wire269)) ^~ forvar283[(1'h0):(1'h0)])) >>> $signed(((!$signed(wire270)) > (-$unsigned(reg273))))))
            begin
              reg285 = $signed($unsigned((((reg280 || forvar278) - (reg282 == (8'hbd))) ?
                  (reg274[(4'he):(4'h8)] ?
                      (wire268 ?
                          (8'hb0) : reg279) : (8'hbb)) : $signed($unsigned(forvar276)))));
              reg286 = ($unsigned(reg277) >>> $signed((((wire268 <<< reg280) ?
                  forvar283 : wire266) * $signed($unsigned(reg273)))));
              reg287 <= (("z" ?
                      $unsigned(wire266) : ($unsigned(forvar283) >= "hqADmm")) ?
                  reg272[(3'h7):(3'h6)] : ((reg274 >>> ((forvar278 <= reg280) ?
                      reg274[(4'he):(3'h4)] : (reg279 ?
                          wire270 : wire269))) >> reg284[(4'h9):(4'h8)]));
              reg288 <= $unsigned($unsigned(reg285[(1'h0):(1'h0)]));
            end
          else
            begin
              reg285 = (~|reg277[(4'ha):(2'h2)]);
              reg286 <= forvar271;
            end
          reg289 <= (8'ha2);
          for (forvar290 = (1'h0); (forvar290 < (2'h2)); forvar290 = (forvar290 + (1'h1)))
            begin
              reg291 <= $signed($unsigned(reg282[(4'h8):(3'h5)]));
              reg292 = (({forvar283,
                      reg280[(2'h2):(2'h2)]} <<< {{(~|(7'h42))}}) ?
                  wire268 : $signed((~reg287)));
            end
          if ($unsigned((-(((8'hae) << (^wire267)) - {(reg272 ?
                  reg291 : forvar271)}))))
            begin
              reg293 <= forvar290;
              reg294 <= reg285[(1'h0):(1'h0)];
            end
          else
            begin
              reg293 <= (8'hb0);
              reg294 = ((^~reg281[(4'hb):(2'h3)]) ?
                  $unsigned((reg288 ?
                      {((8'ha1) | (7'h40))} : reg284[(4'h9):(2'h2)])) : $unsigned($unsigned((~&wire266[(2'h3):(2'h2)]))));
            end
        end
      reg295 = reg288[(4'hf):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg296 = $unsigned($unsigned((reg277 ?
          (~^$unsigned(reg275)) : $signed(reg286))));
      for (forvar297 = (1'h0); (forvar297 < (1'h1)); forvar297 = (forvar297 + (1'h1)))
        begin
          if ((8'had))
            begin
              reg298 = (+($signed(reg288[(2'h2):(1'h1)]) ?
                  (((8'h9f) | (forvar290 ?
                      reg275 : wire265)) || ($signed(forvar276) ~^ reg289)) : ($unsigned($unsigned(reg287)) - forvar297[(3'h5):(3'h5)])));
              reg299 <= (forvar290[(4'h8):(2'h2)] - reg274);
              reg300 <= ($unsigned(($signed((~^forvar297)) >= {(|forvar271)})) ?
                  $signed(reg298[(5'h10):(2'h2)]) : $signed({wire266}));
              reg301 = reg285[(2'h2):(1'h1)];
            end
          else
            begin
              reg298 <= $signed(reg273);
              reg299 <= $unsigned({$signed(forvar290[(4'hd):(4'ha)]),
                  reg281[(4'h8):(3'h7)]});
              reg300 <= $signed((~&forvar283));
              reg301 = $unsigned(reg289);
            end
          reg302 = $signed($unsigned({{(reg301 == reg291)},
              ({(8'haa)} == forvar278[(5'h11):(1'h0)])}));
          reg303 <= reg289[(1'h1):(1'h0)];
        end
      if ((!$signed($unsigned(forvar297))))
        begin
          reg304 = (($unsigned(({reg288, (8'had)} ?
                  reg303 : forvar297[(1'h0):(1'h0)])) || $unsigned($unsigned(reg280[(1'h0):(1'h0)]))) ?
              $unsigned((+(^~(reg287 <= wire268)))) : $unsigned((+reg299[(2'h2):(2'h2)])));
          if (forvar290)
            begin
              reg305 <= (forvar290 >> (wire267 > (|$signed((~forvar276)))));
              reg306 <= (({forvar283, $unsigned($unsigned(reg285))} > (8'h9f)) ?
                  (8'hb5) : reg274);
              reg307 <= (-reg272);
              reg308 <= forvar276[(3'h6):(3'h4)];
              reg309 = reg275[(3'h4):(1'h1)];
            end
          else
            begin
              reg305 <= $unsigned($signed($unsigned((&forvar290[(1'h0):(1'h0)]))));
            end
          if ($unsigned((&(reg303[(5'h15):(5'h11)] ? (-reg279) : reg308))))
            begin
              reg310 <= "CqzRy95";
            end
          else
            begin
              reg310 <= $signed(((-($signed(forvar283) ?
                  wire269[(3'h7):(3'h7)] : reg293[(5'h10):(3'h6)])) <<< {(~|$signed(reg299))}));
              reg311 = ((~^reg272) ?
                  $unsigned(reg284) : $unsigned(((~"Xdqk3no1AmFIC9Lrw") ?
                      {(wire269 < forvar283),
                          "ELUc5b475hWZs1MDPN"} : {(|reg294)})));
              reg312 = ($unsigned($unsigned(((forvar297 & reg300) ?
                  reg273[(3'h7):(3'h4)] : (reg280 << reg291)))) & $signed((^$signed(forvar271))));
              reg313 = {($signed((wire270 ?
                      reg287[(4'hd):(3'h6)] : {(8'hb5),
                          reg275})) < {$unsigned(((8'hb9) ?
                          forvar271 : (7'h43))),
                      reg305[(3'h7):(3'h5)]}),
                  ($unsigned((-$signed((8'hb0)))) ?
                      (^~reg307[(3'h4):(2'h3)]) : reg312)};
              reg314 = $signed(forvar283);
            end
        end
      else
        begin
          reg304 <= reg304[(1'h0):(1'h0)];
          if ((forvar276 ?
              $unsigned((((reg273 ? reg287 : (8'ha3)) > reg288[(1'h0):(1'h0)]) ?
                  reg288[(1'h0):(1'h0)] : reg279)) : $signed((8'hab))))
            begin
              reg305 <= $unsigned(reg296[(4'hc):(4'hc)]);
              reg306 <= reg286[(3'h5):(3'h4)];
              reg307 <= ((forvar283[(2'h2):(2'h2)] ?
                  (^reg313[(4'hc):(4'h8)]) : $unsigned("v19")) ~^ ((((&forvar290) ?
                          (reg277 == reg287) : $signed((8'ha0))) ?
                      ((8'hbc) ?
                          $unsigned(reg277) : $unsigned(reg296)) : ($unsigned(reg277) << reg314)) ?
                  $unsigned(($unsigned(reg304) ?
                      (^reg293) : (reg300 * reg292))) : "B9IglbK3q"));
              reg308 <= (~(($unsigned(wire270) || reg311[(1'h1):(1'h1)]) ?
                  {((reg285 != reg292) ? (^reg308) : {reg281, reg291}),
                      (~^reg296[(4'ha):(3'h5)])} : forvar276));
            end
          else
            begin
              reg305 <= (~|(+$signed($unsigned((reg293 <<< reg288)))));
              reg306 = reg293[(3'h7):(3'h7)];
              reg307 = reg302;
              reg308 <= (7'h40);
              reg309 <= reg279[(1'h1):(1'h0)];
            end
          if ($unsigned(((((reg275 & reg299) ?
                  $signed(reg308) : (8'ha0)) <<< $unsigned($unsigned((8'ha9)))) ?
              $signed($signed({wire270})) : {$signed(reg274[(3'h7):(1'h0)])})))
            begin
              reg310 <= forvar271;
              reg311 <= reg284[(1'h1):(1'h0)];
              reg312 = ((~^$signed(((&(8'hb5)) != (forvar297 ?
                      forvar271 : (8'hbd))))) ?
                  reg300 : ($signed(reg286) + $signed($unsigned($unsigned((8'hbd))))));
              reg313 <= reg307[(3'h4):(2'h2)];
              reg314 <= (+(7'h41));
            end
          else
            begin
              reg310 = (+reg301[(5'h10):(2'h2)]);
              reg311 = $unsigned(reg277[(4'hc):(3'h6)]);
            end
          for (forvar315 = (1'h0); (forvar315 < (1'h0)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 = $unsigned($unsigned($signed(reg304[(2'h3):(1'h1)])));
            end
        end
      if ($unsigned(wire269))
        begin
          if (reg296[(2'h3):(2'h2)])
            begin
              reg317 <= $signed(({($signed(reg299) <= (&reg274)), reg305} ?
                  (~(~&forvar290)) : (((^reg281) || $signed(reg299)) <<< (&$signed((7'h41))))));
              reg318 = (^$signed((~&$signed("18TSrqLBxbfUqZu"))));
              reg319 = $signed((|$signed($unsigned({reg282, reg292}))));
              reg320 = (&$signed(((reg299 != (8'hb5)) ?
                  (&(!reg281)) : reg304[(2'h2):(2'h2)])));
              reg321 = $unsigned(($signed(reg295) ?
                  "l0G9G4Orc6B6kXR6" : $signed(reg306[(4'h9):(2'h2)])));
            end
          else
            begin
              reg317 = $unsigned($signed($unsigned(reg284)));
            end
          if ((({reg279[(4'h8):(4'h8)]} ?
              reg307[(3'h6):(1'h0)] : (reg301 ?
                  $signed($signed(wire267)) : {(-(8'hac))})) | {{$unsigned(((8'h9d) ?
                      (8'ha2) : reg320)),
                  reg277},
              reg272}))
            begin
              reg322 <= ({reg312[(3'h6):(2'h2)]} ?
                  ($signed(({forvar315} ?
                      reg291[(4'hb):(3'h7)] : $unsigned(forvar278))) & $signed({wire265[(1'h1):(1'h1)]})) : (~&(reg273[(2'h3):(2'h2)] == (+reg277[(4'h8):(3'h7)]))));
              reg323 <= ($unsigned("k2dynWlSTi0y57EtSv") ?
                  $unsigned(($signed((reg279 && forvar278)) + (!(~&reg288)))) : reg291);
              reg324 <= wire270;
              reg325 <= ($signed(reg302) ?
                  $signed(((7'h44) * reg281)) : $unsigned({$signed($signed((8'hae))),
                      $signed($signed((8'hac)))}));
            end
          else
            begin
              reg322 <= (&{($unsigned({reg287}) ?
                      ($unsigned(reg325) ?
                          $signed(reg295) : ((8'ha7) ?
                              (8'hbb) : (8'hbc))) : ((^~(8'hae)) ?
                          {reg295, (8'hbb)} : $signed(wire268)))});
              reg323 = $unsigned(($unsigned(($unsigned(reg296) != $unsigned(forvar278))) ?
                  reg311[(1'h0):(1'h0)] : (7'h44)));
              reg324 = reg303[(3'h6):(3'h4)];
              reg325 <= {reg317[(2'h2):(1'h1)],
                  ((((8'ha4) ? ((8'hbc) ? reg281 : reg308) : {forvar315}) ?
                      reg299 : wire266) - $signed(reg300[(3'h5):(3'h5)]))};
            end
        end
      else
        begin
          for (forvar317 = (1'h0); (forvar317 < (1'h0)); forvar317 = (forvar317 + (1'h1)))
            begin
              reg318 <= $signed((|(reg281 + reg286)));
              reg319 <= ((-{(^reg284)}) ?
                  ((8'ha9) ?
                      forvar283[(1'h0):(1'h0)] : $unsigned({(8'hab)})) : reg312);
            end
          for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
            begin
              reg321 = ($unsigned((~|reg291)) - forvar271[(1'h0):(1'h0)]);
              reg322 = ($unsigned(((8'ha0) >> reg281)) ?
                  $unsigned((|((reg279 ? reg285 : reg284) ?
                      (&(8'hbb)) : (forvar320 ?
                          reg301 : (8'hae))))) : (^~(((reg300 <= forvar297) ?
                          $signed(reg317) : (~&reg313)) ?
                      ((~(8'ha4)) ?
                          (!reg291) : reg272[(4'h8):(3'h4)]) : (reg322[(3'h6):(3'h5)] ^ (reg287 << forvar290)))));
              reg323 <= ((((!(reg288 - reg304)) < ($signed(reg302) | reg305)) ^ {(+(reg304 > reg320)),
                      $signed((8'hac))}) ?
                  {(wire267 ? "3VM1gtyGbn3GSEMLp" : "")} : (8'hb7));
              reg324 = (forvar278 << $signed(reg316));
              reg325 <= ({(-{(^~reg323), (-(8'hac))}), (-reg289)} ?
                  $unsigned((-$signed($signed(reg293)))) : {"lz"});
            end
          reg326 = ((reg287 ?
              wire268[(2'h2):(1'h0)] : $signed($signed("aBozz69qLcpDTNXU"))) && reg300[(2'h2):(1'h1)]);
        end
    end
  assign wire327 = forvar297[(4'hc):(3'h4)];
  always
    @(posedge clk) begin
      reg328 <= (({forvar283, ((wire268 ? reg320 : wire268) <= {(8'hb3)})} ?
              {(~&(&forvar271))} : reg314[(5'h10):(5'h10)]) ?
          $signed(reg300[(2'h3):(1'h0)]) : reg307[(2'h2):(2'h2)]);
      reg329 <= (~^($unsigned(((-reg284) >>> (reg307 * reg272))) - $unsigned(((8'hbf) <<< ((8'ha4) & (8'hb2))))));
      for (forvar330 = (1'h0); (forvar330 < (2'h2)); forvar330 = (forvar330 + (1'h1)))
        begin
          for (forvar331 = (1'h0); (forvar331 < (2'h3)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 = reg273[(3'h5):(1'h0)];
              reg333 = (reg305 ?
                  ((~|$signed(wire265)) ?
                      $unsigned((&reg296)) : (~$signed((|reg294)))) : reg319);
              reg334 <= wire266;
            end
          reg335 = $unsigned((^$signed(reg312[(1'h1):(1'h1)])));
          if (reg277[(3'h5):(1'h1)])
            begin
              reg336 <= ($signed((((reg334 >= (8'h9d)) == $signed(reg296)) ?
                      wire270 : (reg286 >> forvar331))) ?
                  ($signed(reg313[(4'hf):(2'h3)]) <= $signed((+reg292[(1'h0):(1'h0)]))) : {(+(^~"rqVRv3Nt5rylh1"))});
              reg337 <= {{$signed((+forvar278[(3'h6):(2'h3)])),
                      (~^(^$signed(wire270)))},
                  reg316[(2'h2):(1'h1)]};
            end
          else
            begin
              reg336 = ($signed((({reg285} <= $signed(reg273)) ?
                      $unsigned($signed(reg328)) : ((reg328 ?
                              reg318 : (8'hbc)) ?
                          $unsigned(reg317) : "A2ogzQN6MYkcn9MVe"))) ?
                  (((8'hb7) | "G") ?
                      $unsigned(reg291[(4'hc):(3'h4)]) : (7'h42)) : $unsigned($unsigned(($signed(forvar315) | $signed(reg323)))));
              reg337 = forvar320[(3'h7):(3'h5)];
              reg338 <= reg310[(1'h1):(1'h0)];
            end
        end
    end
  assign wire339 = reg334;
  always
    @(posedge clk) begin
      for (forvar340 = (1'h0); (forvar340 < (1'h1)); forvar340 = (forvar340 + (1'h1)))
        begin
          for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 = (8'hb3);
              reg343 = reg292;
              reg344 = $signed({(~$signed((-forvar320)))});
            end
          for (forvar345 = (1'h0); (forvar345 < (2'h2)); forvar345 = (forvar345 + (1'h1)))
            begin
              reg346 = (+forvar290);
              reg347 <= (reg310[(3'h5):(3'h4)] <= reg317);
              reg348 <= $signed(reg277);
            end
          reg349 = $signed(forvar276[(2'h2):(2'h2)]);
          reg350 = ({$signed(($unsigned(reg328) <= (^~(8'hb2))))} ?
              ($unsigned(reg279[(2'h2):(1'h1)]) >>> {(|(^(8'haf))),
                  ($signed(reg323) ~^ {wire269})}) : (({$unsigned((8'ha1)),
                          (!reg306)} ?
                      (~^$signed(reg302)) : ({reg346, (8'ha2)} ?
                          (reg288 >= forvar315) : (~|reg285))) ?
                  ($unsigned({reg329,
                      (8'hae)}) & ((~^wire327) ^ wire265[(3'h5):(2'h2)])) : $signed((!{reg326,
                      forvar320}))));
        end
      for (forvar351 = (1'h0); (forvar351 < (2'h2)); forvar351 = (forvar351 + (1'h1)))
        begin
          for (forvar352 = (1'h0); (forvar352 < (1'h0)); forvar352 = (forvar352 + (1'h1)))
            begin
              reg353 <= (~&((~(reg294[(3'h4):(1'h1)] ?
                      (wire267 ? reg282 : reg279) : reg296)) ?
                  $signed(wire267) : forvar352));
              reg354 <= (reg304 ? (8'hb7) : {reg318});
              reg355 = (7'h44);
            end
          reg356 <= (reg324[(2'h2):(1'h0)] * {($signed((reg348 - reg334)) ?
                  (+(+reg302)) : forvar340[(4'h9):(3'h7)]),
              ((reg337 >= ((8'hbe) ?
                  wire265 : (8'hb4))) & $signed((|forvar317)))});
          for (forvar357 = (1'h0); (forvar357 < (1'h0)); forvar357 = (forvar357 + (1'h1)))
            begin
              reg358 = (+reg336[(1'h0):(1'h0)]);
              reg359 <= $signed((~|$signed(((wire269 ?
                  wire265 : wire266) >> reg329))));
              reg360 <= reg335;
              reg361 <= ("gcww14S" ?
                  {((reg307[(4'ha):(2'h3)] ?
                              (wire327 != reg296) : (forvar352 <= reg272)) ?
                          $signed(reg303[(3'h4):(1'h1)]) : ($signed(reg294) | (reg348 ~^ reg307))),
                      reg293[(2'h3):(2'h2)]} : (!$signed(({reg334,
                      forvar317} ^ reg333))));
              reg362 = (~|(reg358[(3'h6):(3'h4)] ?
                  (forvar331 ?
                      $signed((-reg318)) : reg318[(2'h3):(1'h1)]) : $unsigned(($signed((8'ha1)) == reg349[(1'h1):(1'h1)]))));
            end
        end
      reg363 <= $unsigned((!("PACNMAbh" - reg286)));
    end
  assign wire364 = $signed(wire265[(3'h4):(2'h2)]);
  assign wire365 = $signed($signed((($unsigned((8'h9d)) & (forvar340 ?
                       forvar331 : reg346)) || reg361)));
  always
    @(posedge clk) begin
      for (forvar366 = (1'h0); (forvar366 < (3'h4)); forvar366 = (forvar366 + (1'h1)))
        begin
          for (forvar367 = (1'h0); (forvar367 < (1'h0)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 = (^~$unsigned(reg308));
              reg369 <= (&$unsigned({((^reg348) ?
                      {reg323, reg279} : reg321[(2'h2):(1'h0)]),
                  {$signed(reg307), ((8'hb4) ? reg285 : wire268)}}));
              reg370 = ((forvar315 | ((^reg316[(5'h11):(5'h10)]) && $signed($unsigned(forvar341)))) ^ $signed(((reg311[(1'h1):(1'h0)] ?
                      $unsigned(reg361) : (reg346 ? forvar345 : reg359)) ?
                  reg344[(3'h7):(3'h7)] : ($signed(forvar330) ?
                      reg361 : $signed(reg279)))));
              reg371 = wire270[(1'h1):(1'h0)];
              reg372 = $signed($signed(($signed((~^forvar352)) ?
                  ($signed(reg295) ?
                      $unsigned(reg338) : $unsigned(reg369)) : (~(^~reg294)))));
            end
          reg373 = reg302[(3'h5):(2'h3)];
        end
      if (((forvar330[(4'hc):(3'h4)] != (($signed(reg310) ?
              $unsigned(reg358) : $signed(reg359)) ?
          reg373 : (!forvar366))) * reg281))
        begin
          reg374 <= ($unsigned($signed($unsigned(reg298))) ?
              wire265 : (|reg304[(1'h0):(1'h0)]));
          for (forvar375 = (1'h0); (forvar375 < (1'h1)); forvar375 = (forvar375 + (1'h1)))
            begin
              reg376 <= (8'h9d);
              reg377 <= (reg333 ?
                  forvar315 : $unsigned(($signed(reg301[(5'h14):(5'h13)]) + reg337[(1'h0):(1'h0)])));
              reg378 <= $signed($unsigned(reg362));
            end
          for (forvar379 = (1'h0); (forvar379 < (3'h4)); forvar379 = (forvar379 + (1'h1)))
            begin
              reg380 = (reg293[(4'h9):(1'h1)] ?
                  forvar375 : $unsigned({reg329[(1'h0):(1'h0)],
                      $signed((reg358 <<< reg369))}));
              reg381 <= $unsigned(reg282);
              reg382 <= reg360[(1'h1):(1'h0)];
              reg383 = forvar330;
              reg384 <= reg322[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg374 <= {reg324};
        end
      for (forvar385 = (1'h0); (forvar385 < (2'h2)); forvar385 = (forvar385 + (1'h1)))
        begin
          for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 <= forvar385[(1'h1):(1'h1)];
              reg388 <= {(~&reg369)};
              reg389 <= (reg374[(1'h0):(1'h0)] < reg312);
              reg390 = $signed($signed($unsigned(((8'h9d) ?
                  {reg289, reg359} : (reg387 && reg353)))));
              reg391 <= (~|reg348[(1'h0):(1'h0)]);
            end
          for (forvar392 = (1'h0); (forvar392 < (3'h4)); forvar392 = (forvar392 + (1'h1)))
            begin
              reg393 <= reg380;
              reg394 <= (^~{(reg306[(4'hc):(4'hb)] + reg374[(4'hb):(3'h6)]),
                  $unsigned("8FkvUPVCiV")});
              reg395 <= (($unsigned({(reg370 >= forvar340),
                          reg378[(3'h5):(1'h0)]}) ?
                      "5xZiqsDnQ2AHAk8k59b2" : forvar283[(1'h0):(1'h0)]) ?
                  ((((~|(8'hb0)) != $unsigned(reg282)) != $unsigned((8'hbb))) ?
                      (~^forvar367) : $signed(reg363[(2'h2):(2'h2)])) : (7'h40));
            end
          for (forvar396 = (1'h0); (forvar396 < (2'h2)); forvar396 = (forvar396 + (1'h1)))
            begin
              reg397 <= reg322;
              reg398 = $unsigned($unsigned(($unsigned($signed(reg286)) ?
                  reg376[(3'h4):(2'h3)] : (^$signed((8'hb2))))));
              reg399 = $unsigned({((((7'h41) < reg356) ?
                      (wire265 & reg303) : {reg295,
                          (8'hb4)}) <<< (|reg285[(1'h1):(1'h0)])),
                  reg334[(4'h8):(4'h8)]});
              reg400 <= (reg383 >= {$unsigned("zO")});
            end
          reg401 <= (^forvar278);
          reg402 <= ((reg362[(4'h9):(3'h7)] == ((&(reg302 ?
              reg285 : reg291)) <= ((reg333 ? forvar379 : reg306) << {reg273,
              reg371}))) <<< (8'ha5));
        end
      reg403 <= $unsigned(($unsigned($signed(reg294)) ?
          ((^reg293[(4'he):(4'hd)]) ?
              {(forvar345 || reg349)} : $signed((8'h9e))) : reg303));
    end
  assign wire404 = {$unsigned((8'hb9)), ({"M"} * wire267[(3'h7):(3'h7)])};
  assign wire405 = $signed((!reg323));
  always
    @(posedge clk) begin
      reg406 <= reg362;
      reg407 <= (8'ha4);
    end
  always
    @(posedge clk) begin
      for (forvar408 = (1'h0); (forvar408 < (3'h4)); forvar408 = (forvar408 + (1'h1)))
        begin
          for (forvar409 = (1'h0); (forvar409 < (1'h1)); forvar409 = (forvar409 + (1'h1)))
            begin
              reg410 = $signed(reg348[(1'h0):(1'h0)]);
              reg411 <= (forvar379[(2'h2):(1'h1)] != "w12Rpv");
              reg412 <= $unsigned((&(^~(reg343[(2'h2):(1'h0)] ?
                  (~&reg277) : reg318))));
              reg413 = (8'ha0);
              reg414 = forvar320;
            end
          reg415 = (reg305[(4'hd):(3'h4)] * (-$signed($signed((reg308 ?
              (8'hae) : reg281)))));
          for (forvar416 = (1'h0); (forvar416 < (3'h4)); forvar416 = (forvar416 + (1'h1)))
            begin
              reg417 <= ({$unsigned($unsigned((+reg342))), forvar317} ?
                  reg414[(3'h7):(3'h7)] : {($signed(forvar297) >> ("Qh" ?
                          ((8'hab) ? (8'ha1) : (8'hac)) : reg274))});
            end
          reg418 <= forvar315[(4'h8):(4'h8)];
        end
      for (forvar419 = (1'h0); (forvar419 < (2'h2)); forvar419 = (forvar419 + (1'h1)))
        begin
          reg420 = reg371;
          reg421 <= (({($unsigned(reg336) | (reg294 ? reg384 : reg323)),
                  ((reg292 ? reg356 : reg353) & (reg368 << forvar396))} ?
              (wire405 ?
                  (reg287[(5'h12):(4'hb)] ?
                      $unsigned((8'ha6)) : (-reg272)) : reg332[(1'h0):(1'h0)]) : $signed((!(~|reg377)))) < ($signed(forvar320[(5'h12):(4'hc)]) <= $unsigned(((8'ha3) ?
              (reg304 <<< reg368) : (forvar340 ? reg282 : reg300)))));
          if ((reg418[(5'h12):(4'h9)] <<< "8cWLf9hN7Fds"))
            begin
              reg422 <= forvar351;
              reg423 <= (|reg370[(2'h2):(1'h1)]);
            end
          else
            begin
              reg422 = reg381[(2'h2):(2'h2)];
              reg423 <= (|$signed($signed(((~&reg368) ?
                  reg411[(4'h9):(3'h4)] : $unsigned(reg407)))));
              reg424 <= (~^(8'hb5));
              reg425 <= $signed((8'hb8));
            end
          for (forvar426 = (1'h0); (forvar426 < (2'h2)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 <= ("rsIttRro7VXqTEp3QMBD" * $signed(reg395));
              reg428 <= (reg359 || (reg333 && reg335[(3'h5):(2'h3)]));
              reg429 <= (((-(!$unsigned((7'h41)))) ?
                      reg322 : (~^{(~|reg338)})) ?
                  $signed(({(|reg363), (reg418 | reg277)} ?
                      {(-(8'ha0))} : $signed(reg373))) : "bzAeoIfIuP");
              reg430 <= $signed($signed($unsigned(forvar396)));
            end
        end
      reg431 = $unsigned((~|"HTOmeFpOL8mNu"));
      for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
        begin
          for (forvar433 = (1'h0); (forvar433 < (2'h3)); forvar433 = (forvar433 + (1'h1)))
            begin
              reg434 <= ($unsigned(reg291) < reg372);
            end
          for (forvar435 = (1'h0); (forvar435 < (3'h4)); forvar435 = (forvar435 + (1'h1)))
            begin
              reg436 <= {"8laKASR3VB2oaQd",
                  ($unsigned((|$signed(reg356))) >= (8'ha2))};
              reg437 <= reg418[(5'h11):(4'hd)];
              reg438 = $signed((reg376 ?
                  ((reg329[(4'ha):(1'h1)] ?
                      $unsigned(reg287) : ((8'hb3) ~^ reg369)) <= $signed((^~reg353))) : (reg321[(1'h1):(1'h1)] >> "kJwOGWF")));
              reg439 <= forvar278;
            end
          if (reg329)
            begin
              reg440 <= {(8'hb5), $signed(forvar320)};
              reg441 = ($unsigned(((reg381[(2'h3):(2'h3)] >> (~&(8'haf))) ?
                  $unsigned($unsigned(reg306)) : (forvar276 << (reg313 ?
                      wire339 : (8'hac))))) > (~{$signed((reg359 ?
                      (8'hb9) : (8'hba)))}));
            end
          else
            begin
              reg440 = reg403;
              reg441 <= ($signed(reg313[(3'h5):(1'h0)]) ?
                  ((((|forvar341) > $unsigned(reg371)) ?
                      ($unsigned(reg427) ?
                          ((8'ha4) * reg406) : "7QXBbP8w") : (!reg440)) < $signed({(~|wire268)})) : reg373[(3'h4):(2'h3)]);
              reg442 <= ($unsigned((($signed(forvar315) || $unsigned(reg295)) ?
                      reg336 : "gMeVgfkiN02ok")) ?
                  "3M371BPwqJ" : $signed(reg292[(1'h1):(1'h1)]));
            end
          for (forvar443 = (1'h0); (forvar443 < (2'h3)); forvar443 = (forvar443 + (1'h1)))
            begin
              reg444 <= {reg391, $signed((8'hb8))};
              reg445 <= (reg319[(4'h9):(1'h1)] ?
                  ($signed($signed($unsigned(reg399))) ?
                      reg343[(1'h1):(1'h0)] : reg387) : (reg322[(2'h2):(2'h2)] ?
                      (reg378[(3'h7):(3'h4)] ?
                          $signed($signed((8'hb4))) : {(|wire268),
                              reg293}) : $unsigned((~|$unsigned(reg349)))));
              reg446 <= {$signed(reg314[(3'h6):(1'h0)])};
              reg447 = $signed((&{reg320[(3'h5):(3'h5)]}));
              reg448 = forvar271[(1'h0):(1'h0)];
            end
        end
      for (forvar449 = (1'h0); (forvar449 < (1'h1)); forvar449 = (forvar449 + (1'h1)))
        begin
          reg450 <= (reg285[(1'h0):(1'h0)] ?
              (reg429[(2'h3):(2'h3)] ? forvar366 : reg350) : reg335);
          for (forvar451 = (1'h0); (forvar451 < (2'h2)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 = ((reg447[(1'h1):(1'h1)] ~^ (reg428[(1'h1):(1'h1)] ?
                  (^~reg280) : reg287[(5'h13):(2'h2)])) << $unsigned(forvar330[(4'h9):(1'h0)]));
              reg453 <= forvar409[(1'h0):(1'h0)];
              reg454 = reg329;
            end
          for (forvar455 = (1'h0); (forvar455 < (2'h3)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 <= (($unsigned($unsigned($unsigned(reg287))) << (forvar367[(4'h8):(4'h8)] | (~|(|reg382)))) <<< ((((reg356 <= reg394) << $signed(reg308)) ?
                  {(reg354 | forvar351),
                      reg344[(4'h9):(1'h1)]} : (&$unsigned(reg440))) * ((&{(8'ha8)}) ?
                  $signed(reg301) : "F7VP")));
              reg457 <= reg415;
              reg458 = ((forvar290[(4'hd):(2'h2)] ~^ reg314[(5'h12):(2'h2)]) - reg444);
              reg459 = $signed((forvar278 ?
                  $unsigned((wire365 | forvar340[(4'ha):(2'h2)])) : (reg401[(2'h2):(2'h2)] <= forvar315)));
            end
          reg460 <= ((&$signed((~(|reg337)))) ^ forvar386[(4'h9):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      if (reg401[(2'h2):(1'h1)])
        begin
          for (forvar461 = (1'h0); (forvar461 < (1'h1)); forvar461 = (forvar461 + (1'h1)))
            begin
              reg462 <= $signed(reg311[(2'h2):(1'h0)]);
              reg463 = $unsigned(reg440);
              reg464 <= reg355;
              reg465 <= ({wire269} == reg417[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          if ((reg384 & $unsigned(((~|(forvar366 ? reg389 : reg427)) ?
              ((reg371 ?
                  (8'ha2) : reg346) ^ (reg400 != reg423)) : ($signed(forvar315) ?
                  reg285[(2'h2):(2'h2)] : reg335[(5'h12):(4'he)])))))
            begin
              reg461 <= $signed($unsigned((($unsigned(forvar433) ?
                      reg369 : ((8'h9e) ? reg313 : reg336)) ?
                  ((reg442 || reg430) ?
                      $unsigned(wire404) : "g7ob3Gm9qonWy2CM") : ($unsigned(wire269) * reg384[(4'hd):(2'h2)]))));
              reg462 = reg442[(4'h9):(2'h2)];
            end
          else
            begin
              reg461 = reg307;
              reg462 = forvar330;
              reg463 = reg328;
              reg464 = $unsigned($signed({((reg332 != reg398) * {reg407,
                      (8'hb8)}),
                  ((8'hb2) || $unsigned(reg387))}));
            end
          reg465 <= forvar290;
          for (forvar466 = (1'h0); (forvar466 < (2'h2)); forvar466 = (forvar466 + (1'h1)))
            begin
              reg467 = (reg291[(4'he):(3'h4)] <<< $unsigned($signed(forvar443)));
              reg468 <= $unsigned(reg281);
              reg469 <= (+({($unsigned(reg323) ?
                          $unsigned(reg338) : (~^reg332)),
                      $signed(reg420)} ?
                  reg295[(4'he):(3'h5)] : ($signed((&reg450)) ^~ (reg401 ?
                      {reg383} : reg380[(5'h11):(4'h9)]))));
              reg470 = "WR45W";
              reg471 = ((reg346 >> (|$unsigned(reg458[(4'h8):(3'h5)]))) ?
                  {reg439} : ((wire270 ?
                          (!(|forvar317)) : $signed($unsigned(reg420))) ?
                      ((-(reg463 ^~ forvar290)) + $unsigned($signed(reg421))) : $signed(($signed(reg442) ^ $signed(wire267)))));
            end
          if ($unsigned(({($unsigned(reg301) ^~ (reg289 <<< reg464)),
              $signed({(8'h9d)})} << $signed(((reg471 == reg460) < reg277)))))
            begin
              reg472 = (&reg358[(3'h5):(3'h4)]);
              reg473 <= $signed($signed($unsigned(($unsigned(reg444) ?
                  "KIRK" : reg387[(4'h9):(1'h1)]))));
            end
          else
            begin
              reg472 <= (+$signed(((8'hb5) == reg320[(4'h8):(1'h0)])));
            end
          if ((-forvar331))
            begin
              reg474 <= (8'hbe);
              reg475 <= {(~&forvar315[(4'h9):(1'h1)]),
                  (reg423[(3'h4):(2'h2)] + reg361)};
            end
          else
            begin
              reg474 <= "ew93pcNWJ";
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module132
#( parameter param260 = (((^(+{(8'h9c), (8'ha8)})) ? (+{(&(8'hb8)), ((8'ha9) ^ (7'h44))}) : ((((8'ha2) & (8'hb8)) ? {(8'hb2), (8'hb4)} : ((7'h40) <= (8'hac))) ? (((8'ha6) != (8'hbe)) ? ((8'hb5) ? (8'hb1) : (8'ha4)) : (8'hac)) : {(+(8'ha0))})) || {(~|(+((8'h9c) - (8'hb1)))), (~&(((8'hae) <<< (7'h42)) ? (^~(8'hb0)) : {(8'ha4), (8'haa)}))}) )
(y, clk, wire137, wire136, wire135, wire134, wire133);
  output wire [(32'h598):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire137;
  input wire [(4'h8):(1'h0)] wire136;
  input wire [(3'h6):(1'h0)] wire135;
  input wire [(5'h12):(1'h0)] wire134;
  input wire [(5'h15):(1'h0)] wire133;
  wire signed [(4'hb):(1'h0)] wire259;
  wire [(3'h4):(1'h0)] wire258;
  wire signed [(4'hb):(1'h0)] wire257;
  reg signed [(4'h9):(1'h0)] reg256 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg254 = (1'h0);
  reg [(3'h6):(1'h0)] reg253 = (1'h0);
  reg [(3'h5):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg250 = (1'h0);
  reg [(4'hb):(1'h0)] reg249 = (1'h0);
  reg [(4'ha):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar247 = (1'h0);
  reg [(5'h14):(1'h0)] reg246 = (1'h0);
  reg [(4'he):(1'h0)] reg245 = (1'h0);
  reg [(4'hb):(1'h0)] reg244 = (1'h0);
  reg [(4'h9):(1'h0)] forvar243 = (1'h0);
  reg [(4'he):(1'h0)] forvar229 = (1'h0);
  reg [(5'h15):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg241 = (1'h0);
  reg [(3'h6):(1'h0)] reg240 = (1'h0);
  reg [(5'h11):(1'h0)] reg239 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar238 = (1'h0);
  reg [(5'h15):(1'h0)] reg237 = (1'h0);
  reg [(4'hf):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(4'hc):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar231 = (1'h0);
  reg [(4'hc):(1'h0)] reg230 = (1'h0);
  reg [(5'h13):(1'h0)] reg229 = (1'h0);
  reg [(5'h11):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg227 = (1'h0);
  reg [(2'h2):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar225 = (1'h0);
  reg [(5'h12):(1'h0)] reg224 = (1'h0);
  reg [(5'h10):(1'h0)] reg223 = (1'h0);
  reg [(4'hb):(1'h0)] reg222 = (1'h0);
  reg [(2'h2):(1'h0)] reg221 = (1'h0);
  reg [(2'h3):(1'h0)] forvar220 = (1'h0);
  reg [(4'ha):(1'h0)] reg219 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg218 = (1'h0);
  reg [(5'h11):(1'h0)] reg217 = (1'h0);
  reg [(5'h14):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg214 = (1'h0);
  reg [(3'h6):(1'h0)] reg213 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg212 = (1'h0);
  reg [(4'he):(1'h0)] forvar211 = (1'h0);
  reg [(5'h14):(1'h0)] reg210 = (1'h0);
  reg [(3'h5):(1'h0)] forvar209 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg208 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar207 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar203 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar201 = (1'h0);
  reg [(2'h3):(1'h0)] reg203 = (1'h0);
  reg [(4'h9):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg201 = (1'h0);
  reg signed [(4'he):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg199 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg198 = (1'h0);
  reg [(5'h15):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg196 = (1'h0);
  reg [(5'h10):(1'h0)] reg195 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar194 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg193 = (1'h0);
  reg [(4'ha):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar191 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg190 = (1'h0);
  reg [(4'hd):(1'h0)] reg189 = (1'h0);
  reg [(3'h4):(1'h0)] reg188 = (1'h0);
  reg [(3'h4):(1'h0)] reg187 = (1'h0);
  reg [(4'hd):(1'h0)] reg186 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg185 = (1'h0);
  reg [(5'h10):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg182 = (1'h0);
  reg [(3'h4):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg180 = (1'h0);
  reg [(3'h4):(1'h0)] forvar179 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar178 = (1'h0);
  reg [(4'ha):(1'h0)] reg177 = (1'h0);
  wire [(4'ha):(1'h0)] wire176;
  reg signed [(3'h7):(1'h0)] reg175 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg173 = (1'h0);
  reg [(3'h4):(1'h0)] reg172 = (1'h0);
  reg [(2'h2):(1'h0)] reg171 = (1'h0);
  reg [(3'h5):(1'h0)] reg168 = (1'h0);
  reg [(4'hc):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg169 = (1'h0);
  reg [(4'he):(1'h0)] forvar168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar166 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg165 = (1'h0);
  reg [(4'h9):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg163 = (1'h0);
  reg [(2'h3):(1'h0)] forvar162 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg161 = (1'h0);
  reg [(3'h5):(1'h0)] reg160 = (1'h0);
  reg [(5'h13):(1'h0)] reg159 = (1'h0);
  reg [(5'h15):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg152 = (1'h0);
  reg [(4'hc):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg149 = (1'h0);
  reg [(5'h14):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg146 = (1'h0);
  reg [(5'h11):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg143 = (1'h0);
  reg [(5'h13):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar141 = (1'h0);
  reg [(4'hd):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg139 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire138;
  assign y = {wire259,
                 wire258,
                 wire257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 forvar247,
                 reg246,
                 reg245,
                 reg244,
                 forvar243,
                 forvar229,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 forvar238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 forvar231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 forvar225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 forvar220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 forvar211,
                 reg210,
                 forvar209,
                 reg208,
                 forvar207,
                 reg206,
                 reg205,
                 reg204,
                 forvar203,
                 forvar201,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 forvar194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 forvar179,
                 forvar178,
                 reg177,
                 wire176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg168,
                 reg166,
                 reg170,
                 reg169,
                 forvar168,
                 reg167,
                 forvar166,
                 reg165,
                 reg164,
                 reg163,
                 forvar162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 forvar157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 forvar151,
                 reg150,
                 reg149,
                 reg148,
                 forvar147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 forvar141,
                 reg140,
                 reg139,
                 wire138,
                 (1'h0)};
  assign wire138 = (^~(~$signed($signed(wire134[(4'ha):(1'h0)]))));
  always
    @(posedge clk) begin
      reg139 = wire133[(4'hd):(2'h2)];
      reg140 <= (($unsigned(($unsigned(wire134) ?
          wire134 : (reg139 ?
              wire137 : wire134))) + (~^((~(8'ha7)) | (8'ha0)))) == $unsigned((($unsigned(wire134) < (8'hb8)) != (~(wire137 * wire133)))));
      for (forvar141 = (1'h0); (forvar141 < (2'h3)); forvar141 = (forvar141 + (1'h1)))
        begin
          if (($signed("tUnmxh") ?
              $unsigned($unsigned(((wire133 ?
                  forvar141 : reg140) == $unsigned(wire134)))) : ($signed(wire133[(4'hc):(2'h3)]) ?
                  ($signed(wire136) <<< (forvar141[(1'h0):(1'h0)] ?
                      wire137[(2'h2):(2'h2)] : "R")) : $signed((8'ha3)))))
            begin
              reg142 = (|$unsigned($signed(((!wire135) ?
                  (!wire138) : wire136))));
              reg143 <= ($signed($signed((!(reg140 - wire137)))) ~^ $signed(($unsigned($unsigned(reg140)) ?
                  wire134[(5'h10):(4'hd)] : $signed((wire134 - reg142)))));
              reg144 <= $unsigned({wire137[(2'h2):(2'h2)]});
            end
          else
            begin
              reg142 <= (^$signed(((^~(+reg142)) ?
                  wire136[(4'h8):(1'h0)] : (wire134 ?
                      $signed(wire133) : reg144))));
              reg143 <= {{((~|(8'ha6)) ?
                          $signed(wire136) : (((8'h9f) ^ wire134) - ((8'hab) ?
                              reg143 : (8'hba)))),
                      wire137},
                  {wire135}};
              reg144 = reg142[(1'h0):(1'h0)];
              reg145 = ((!(((wire137 == forvar141) == reg139[(3'h6):(1'h0)]) ?
                      {reg140[(3'h6):(2'h3)],
                          (&(8'ha0))} : ($unsigned(forvar141) ?
                          (+reg144) : $signed(wire134)))) ?
                  wire135[(1'h1):(1'h1)] : (((reg143 + (^~(8'hb3))) ^~ reg139[(5'h11):(1'h1)]) ?
                      wire138 : reg142[(1'h0):(1'h0)]));
              reg146 = "h9CfW7gUvO5UwUbY2";
            end
          for (forvar147 = (1'h0); (forvar147 < (1'h1)); forvar147 = (forvar147 + (1'h1)))
            begin
              reg148 <= ({$signed((!(reg142 ? reg146 : reg139)))} ?
                  (~&(^~wire137)) : $unsigned($unsigned((|$signed(wire138)))));
              reg149 <= {$unsigned($unsigned(wire135[(1'h0):(1'h0)]))};
            end
          reg150 <= reg145;
          for (forvar151 = (1'h0); (forvar151 < (2'h2)); forvar151 = (forvar151 + (1'h1)))
            begin
              reg152 = wire136;
              reg153 = (-reg152[(1'h1):(1'h1)]);
              reg154 <= $signed(($signed($signed($unsigned(reg152))) ?
                  wire134[(4'he):(3'h6)] : forvar151));
              reg155 <= ($signed(((^~reg149) >= (-((8'hb2) ^~ forvar147)))) & (~&{reg145}));
              reg156 = $signed(($unsigned(reg153) ^~ reg149[(4'h9):(2'h3)]));
            end
          for (forvar157 = (1'h0); (forvar157 < (2'h2)); forvar157 = (forvar157 + (1'h1)))
            begin
              reg158 = $signed($signed($unsigned($signed({wire136, (8'ha2)}))));
              reg159 = ((~^(^$unsigned((~|wire133)))) ?
                  wire136[(1'h1):(1'h1)] : (|((8'ha5) | (~{reg142, reg145}))));
              reg160 <= $unsigned($signed((reg152 ?
                  reg142[(4'he):(3'h4)] : reg159[(2'h3):(2'h2)])));
            end
        end
      reg161 = $signed({reg152, {{wire136[(1'h1):(1'h1)]}}});
    end
  always
    @(posedge clk) begin
      if ($unsigned({(~(((7'h41) || reg150) ?
              (reg149 ? reg152 : reg156) : {reg152, wire137}))}))
        begin
          for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 <= reg144;
              reg164 <= $signed(wire134);
              reg165 = {(reg144 ?
                      ((+(wire135 ?
                          (8'haf) : reg144)) >= $signed((~|reg161))) : (~^reg164[(2'h3):(2'h3)])),
                  $unsigned($unsigned(((wire134 ~^ (8'hb4)) ?
                      (~^reg156) : "reZv1N")))};
            end
          for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 = {wire134};
            end
          for (forvar168 = (1'h0); (forvar168 < (3'h4)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 = $signed(reg149[(4'hb):(3'h4)]);
            end
          reg170 <= $signed({$signed($unsigned($signed(reg148)))});
        end
      else
        begin
          for (forvar162 = (1'h0); (forvar162 < (2'h2)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 <= $unsigned(reg160[(3'h5):(2'h3)]);
              reg164 = reg145;
              reg165 <= reg170;
              reg166 = wire134[(4'hb):(2'h3)];
              reg167 <= (wire133 ^ (-(reg148 > {(reg161 <<< reg139),
                  $unsigned(reg161)})));
            end
          if ((($signed(((8'hbd) << (~&reg169))) ?
                  ((8'ha0) ?
                      ((reg154 << reg154) <= $signed(reg155)) : {((8'hbd) ~^ forvar162),
                          (forvar151 ?
                              (8'hb4) : reg163)}) : ((reg148[(4'hc):(1'h0)] ?
                      (~&reg140) : (wire136 << reg149)) > {$signed(reg146)})) ?
              ($unsigned(({reg158} ? (|(8'ha9)) : $unsigned(forvar157))) ?
                  {forvar141[(1'h0):(1'h0)],
                      reg160[(2'h3):(2'h3)]} : $signed($unsigned({reg152}))) : (~($unsigned((forvar147 ?
                      forvar151 : (8'haa))) ?
                  (8'hb6) : reg152))))
            begin
              reg168 = "STNaUG2xTo60I1HZwQ";
            end
          else
            begin
              reg168 <= (((^~{reg167[(2'h3):(1'h0)]}) & wire138) ?
                  "YOaGcJctfHYAwJFYs" : reg163);
              reg169 <= wire134;
              reg170 = reg167;
              reg171 = (($signed(((|forvar141) ? wire136 : {forvar151})) ?
                  (($signed(reg161) ?
                          (reg156 ? (8'ha2) : (7'h42)) : (+forvar147)) ?
                      forvar147 : $signed($unsigned(reg152))) : reg143) > "dp");
              reg172 <= $signed($signed(forvar141));
            end
          if (($unsigned((~&((^reg153) ? $signed(reg155) : reg160))) ?
              ($signed(reg148) ?
                  ({reg159,
                      $unsigned(wire136)} ^ {forvar162[(1'h1):(1'h1)]}) : $unsigned(forvar151)) : {((reg149 * (-reg166)) - wire138),
                  $signed((reg161[(1'h1):(1'h1)] ?
                      (reg139 ? reg170 : reg166) : reg167))}))
            begin
              reg173 = (!$unsigned(($unsigned($signed(reg149)) >= (^~reg142[(5'h11):(3'h5)]))));
              reg174 <= $unsigned((^reg148));
            end
          else
            begin
              reg173 <= reg144;
            end
          reg175 = $signed($unsigned($signed(forvar141)));
        end
    end
  assign wire176 = $signed(($unsigned(((8'hbd) >= wire137[(2'h2):(1'h0)])) << "aJ9pQRrlIVPGMuzZzp"));
  always
    @(posedge clk) begin
      reg177 <= (~($signed((|reg155[(3'h7):(1'h0)])) + $unsigned((~reg140))));
      for (forvar178 = (1'h0); (forvar178 < (1'h1)); forvar178 = (forvar178 + (1'h1)))
        begin
          for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
            begin
              reg180 = $signed(reg160[(1'h0):(1'h0)]);
              reg181 <= (~|(~|reg144[(3'h7):(3'h7)]));
              reg182 <= ($signed((reg165[(1'h0):(1'h0)] && reg139)) >> $unsigned({$signed("")}));
              reg183 = ({(-{reg159}),
                  ($unsigned({(8'ha2)}) ?
                      (-((8'hb9) != reg170)) : wire135)} << (((&{reg181}) ?
                  $signed((8'ha7)) : (reg152 ?
                      forvar166[(4'hf):(4'he)] : forvar147[(3'h5):(3'h5)])) ~^ (~^{$unsigned(forvar168),
                  reg142})));
              reg184 = ($signed(($signed((wire138 == (8'haf))) ?
                  (reg177[(2'h2):(1'h0)] == (~&reg158)) : $unsigned((8'hb8)))) || forvar141);
            end
          reg185 = (|(((+reg168) ?
                  (reg156 ?
                      (reg152 ?
                          reg168 : forvar157) : wire135[(1'h0):(1'h0)]) : wire133) ?
              ($signed(forvar162) > (wire136 ^~ (forvar166 != forvar162))) : {{$signed(reg152)}}));
          if ($signed($unsigned({{$unsigned((8'haa)), $signed(reg150)},
              (reg145[(4'hf):(3'h6)] & wire176)})))
            begin
              reg186 <= reg158;
              reg187 = reg139;
              reg188 = $unsigned((reg172 - reg183[(3'h6):(1'h1)]));
              reg189 = reg186[(4'hb):(4'hb)];
              reg190 <= $signed({(reg155 ?
                      (^~(|reg165)) : $signed((reg172 == forvar179)))});
            end
          else
            begin
              reg186 <= $unsigned($unsigned($unsigned(forvar166[(4'ha):(2'h2)])));
              reg187 <= (&wire138);
              reg188 <= (|{((~reg180[(1'h0):(1'h0)]) <= ((&wire176) != "qwPMoWsg1U327i"))});
              reg189 <= $unsigned(("92oKRZd6hc3" ? reg187 : reg190));
            end
          for (forvar191 = (1'h0); (forvar191 < (2'h3)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= (^($signed(reg182[(3'h6):(1'h0)]) && (reg150 ?
                  ({forvar151, reg164} ?
                      $unsigned(reg154) : $unsigned(reg175)) : {$unsigned(wire133)})));
              reg193 = {{wire133}};
            end
          for (forvar194 = (1'h0); (forvar194 < (2'h2)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg195 <= (~|$unsigned(reg184[(2'h3):(2'h3)]));
              reg196 <= $signed("toqkG2wNcBti49VtqlK");
            end
        end
      reg197 = reg161;
      reg198 <= {{reg153},
          $unsigned($signed(((8'hba) ?
              (reg153 ? reg193 : reg168) : $unsigned((8'hb7)))))};
      reg199 = $unsigned((8'ha9));
    end
  always
    @(posedge clk) begin
      if ((~forvar147[(3'h4):(1'h0)]))
        begin
          reg200 <= (8'hbb);
          if ((~^(($unsigned((reg182 > reg181)) ?
              $unsigned($signed((8'hb9))) : $signed($unsigned(wire135))) - $unsigned($signed("fWDKFyMoLVvD8Sm27Stc")))))
            begin
              reg201 = forvar166;
              reg202 = $unsigned((^$signed({$signed(reg173)})));
              reg203 = $signed((~((reg153 < (reg189 ^ reg144)) + reg161[(2'h2):(1'h0)])));
            end
          else
            begin
              reg201 = (~^("VCMQA" ?
                  (reg154 ^ $signed(reg143[(3'h4):(2'h2)])) : (-reg160[(3'h4):(1'h0)])));
            end
        end
      else
        begin
          reg200 <= $unsigned((|((reg160 ? (^~reg182) : (reg190 >> (8'had))) ?
              (^~(~reg184)) : forvar194[(1'h1):(1'h1)])));
          for (forvar201 = (1'h0); (forvar201 < (3'h4)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 = $unsigned($signed(reg154));
            end
          for (forvar203 = (1'h0); (forvar203 < (1'h1)); forvar203 = (forvar203 + (1'h1)))
            begin
              reg204 <= (^~{forvar194[(2'h2):(1'h0)], wire137[(1'h0):(1'h0)]});
              reg205 = $unsigned(reg193[(4'he):(4'hb)]);
              reg206 <= {$signed($unsigned($unsigned(reg171[(1'h0):(1'h0)]))),
                  ({forvar166} ?
                      $unsigned((+$unsigned(reg171))) : ((reg204[(1'h0):(1'h0)] ^ forvar157[(2'h2):(1'h0)]) ?
                          $signed((wire135 || reg142)) : forvar151))};
            end
          for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 <= ($signed($signed($unsigned((wire136 ?
                  reg199 : forvar168)))) == reg182);
            end
          for (forvar209 = (1'h0); (forvar209 < (1'h1)); forvar209 = (forvar209 + (1'h1)))
            begin
              reg210 = $unsigned((($unsigned((reg148 & reg156)) ?
                  reg164[(2'h3):(2'h3)] : (~(reg168 ?
                      reg177 : reg199))) ^ forvar201[(4'ha):(4'ha)]));
            end
        end
      for (forvar211 = (1'h0); (forvar211 < (2'h2)); forvar211 = (forvar211 + (1'h1)))
        begin
          if (reg144)
            begin
              reg212 <= $unsigned((^~"QfJohq88i"));
              reg213 <= reg206;
              reg214 <= (|($signed((-(reg173 << forvar178))) ?
                  (^($signed(reg156) ?
                      $unsigned(reg189) : wire133[(1'h1):(1'h1)])) : (&reg149)));
              reg215 <= {(!"MWdlVQ")};
            end
          else
            begin
              reg212 <= reg142;
              reg213 = ($unsigned($unsigned(reg198[(1'h0):(1'h0)])) <= $signed(reg183));
              reg214 = ("Y" ?
                  {{(reg197[(4'ha):(4'h9)] ?
                              reg156 : (reg160 ? reg182 : reg154))},
                      ((7'h44) ?
                          reg200[(4'hc):(3'h6)] : (8'ha6))} : (^~((^~$signed(reg173)) & $unsigned($signed(forvar194)))));
            end
          if ((((&$signed($signed((8'ha1)))) - (reg212[(4'h8):(3'h5)] > (~reg175))) + reg172))
            begin
              reg216 = $unsigned($signed((~^reg190[(1'h0):(1'h0)])));
              reg217 = reg215[(3'h4):(1'h0)];
              reg218 = reg140;
            end
          else
            begin
              reg216 = reg192;
              reg217 <= forvar211;
              reg218 <= reg164[(2'h3):(2'h2)];
              reg219 = (reg216[(4'h9):(4'h9)] <= ((8'ha7) + ({$unsigned(reg150)} ?
                  reg154 : reg154[(1'h0):(1'h0)])));
            end
          for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
            begin
              reg221 <= ($unsigned((&$signed(reg145))) > (~&reg177));
              reg222 <= ((8'hbe) ?
                  wire138 : ($unsigned($unsigned(reg159[(3'h6):(1'h1)])) ?
                      (((~^reg144) && (reg219 <<< (8'hba))) - (^~reg158)) : reg163[(2'h2):(1'h1)]));
            end
          reg223 = reg201;
          reg224 = $signed($unsigned(reg154));
        end
      if ((!reg160[(1'h1):(1'h0)]))
        begin
          for (forvar225 = (1'h0); (forvar225 < (2'h3)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= $unsigned(reg140[(1'h1):(1'h0)]);
              reg227 <= (reg216[(5'h13):(5'h13)] && ((8'hb4) > reg153[(4'ha):(1'h0)]));
              reg228 <= reg223[(2'h2):(1'h1)];
              reg229 = ((((^~$signed((8'hb2))) - ($signed(reg166) < $signed(reg177))) ?
                  {$signed($signed(reg172))} : (((reg173 ?
                      reg175 : (7'h41)) + forvar225[(3'h6):(3'h6)]) || (~|(!(8'ha9))))) && reg160);
              reg230 <= $signed(wire134[(2'h3):(1'h0)]);
            end
          for (forvar231 = (1'h0); (forvar231 < (3'h4)); forvar231 = (forvar231 + (1'h1)))
            begin
              reg232 <= ({reg223[(4'hb):(4'hb)]} ?
                  $unsigned(reg186[(4'ha):(4'h9)]) : ((({(8'hae),
                          reg146} > forvar194) && (|reg190[(4'h9):(3'h7)])) ?
                      (&$unsigned((~|forvar191))) : (+$unsigned(reg195[(4'h8):(3'h4)]))));
              reg233 <= reg213;
              reg234 <= "vrLoYDY";
              reg235 <= $unsigned({($unsigned(reg223[(4'h9):(3'h7)]) ?
                      (reg170 ? wire133 : ((8'hbe) & reg228)) : reg139)});
            end
          reg236 = reg168;
          reg237 = $unsigned((reg172 ^ reg163));
          for (forvar238 = (1'h0); (forvar238 < (2'h3)); forvar238 = (forvar238 + (1'h1)))
            begin
              reg239 <= reg195;
              reg240 <= $signed((~&{""}));
              reg241 <= (^$unsigned((reg228 ?
                  forvar231 : $signed((^(7'h42))))));
              reg242 = (~|($unsigned((reg208[(4'hb):(1'h1)] ?
                  forvar157[(1'h1):(1'h0)] : $signed(reg219))) > $unsigned(((!(8'hb7)) <= forvar162))));
            end
        end
      else
        begin
          for (forvar225 = (1'h0); (forvar225 < (1'h1)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 = $unsigned({(reg210[(4'hf):(3'h6)] ?
                      $signed((reg212 << (8'ha4))) : (^reg165[(2'h2):(1'h1)])),
                  reg144});
              reg227 = (reg159[(4'h8):(2'h2)] ?
                  ((+$signed($unsigned(reg239))) ^~ "bXsuWBy0MNZgF4s9q") : reg159);
              reg228 <= ((!(8'h9d)) ? reg142[(3'h6):(1'h0)] : (!forvar166));
            end
          for (forvar229 = (1'h0); (forvar229 < (2'h2)); forvar229 = (forvar229 + (1'h1)))
            begin
              reg230 = (reg180 ?
                  $signed((((-reg142) ? (|(8'hbc)) : (!(8'ha8))) ?
                      reg181[(1'h0):(1'h0)] : $signed((forvar209 ?
                          reg167 : reg182)))) : $signed(reg224[(4'hb):(2'h3)]));
            end
          for (forvar231 = (1'h0); (forvar231 < (1'h1)); forvar231 = (forvar231 + (1'h1)))
            begin
              reg232 = (8'hb7);
              reg233 = ((($signed((reg182 ^ reg144)) <= {$unsigned(reg169)}) ?
                  wire135[(3'h5):(3'h5)] : ("odSdzDh8LzzWG" || (((8'hbe) ?
                          (8'hbc) : reg228) ?
                      (!reg197) : {(7'h43)}))) ^~ {(|{$signed(forvar162)}),
                  (($signed((8'hba)) > (forvar166 ? wire176 : reg193)) ?
                      ($unsigned((8'ha4)) ?
                          {reg222,
                              reg198} : forvar229[(4'he):(3'h4)]) : $signed((forvar141 ?
                          reg219 : reg218)))});
            end
        end
      if (($unsigned(((((8'hb2) ? reg170 : reg173) ?
              $signed((8'ha7)) : reg240) ?
          (-(~(8'ha1))) : ($unsigned(reg222) ?
              $unsigned((8'hb4)) : $unsigned((8'haf))))) >> reg216[(3'h5):(3'h4)]))
        begin
          for (forvar243 = (1'h0); (forvar243 < (1'h1)); forvar243 = (forvar243 + (1'h1)))
            begin
              reg244 = (|reg144);
              reg245 <= (~&$unsigned(($signed("xEkbpXeMIvbOcXIJZB") ?
                  $unsigned(reg222) : ((|reg215) - $unsigned(reg154)))));
              reg246 <= $unsigned((wire136 ?
                  "Lc9LzcmEICML" : ($unsigned((8'hb7)) ?
                      $signed(reg159[(5'h12):(3'h5)]) : (~&$unsigned(forvar209)))));
            end
          for (forvar247 = (1'h0); (forvar247 < (1'h0)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= reg140;
              reg249 <= ({$unsigned(((wire176 ?
                      reg183 : reg237) && (~reg233)))} > ({forvar168} ?
                  ($unsigned((reg195 >= reg186)) ?
                      (~reg208) : $unsigned((^reg202))) : {(~^(^~reg212)),
                      (^forvar179[(1'h0):(1'h0)])}));
              reg250 = reg180[(4'he):(1'h0)];
              reg251 = reg227;
            end
          if ((reg232[(4'hd):(3'h6)] ?
              {$unsigned($unsigned($signed(reg203)))} : reg216))
            begin
              reg252 = "aDmTR4yPRVexSpW8LH";
              reg253 <= reg252;
              reg254 <= ((+($unsigned(reg183[(4'hc):(3'h7)]) ?
                  ((reg189 * reg187) ^ reg218[(2'h2):(2'h2)]) : (-reg195))) ^~ $unsigned(reg150[(3'h6):(2'h2)]));
              reg255 = forvar151;
            end
          else
            begin
              reg252 <= ($signed(({(wire176 - (8'haf)),
                      {forvar203}} >> $unsigned(reg224[(4'hd):(4'hc)]))) ?
                  $signed({{$unsigned(reg196),
                          ((8'ha0) ~^ forvar238)}}) : $signed((forvar194 - {reg246[(3'h7):(3'h6)]})));
              reg253 <= {(^~(((reg156 ^~ reg144) ?
                          "3MYytzMX1a0ffwqcg" : reg171) ?
                      wire138[(1'h1):(1'h1)] : ((~reg166) ?
                          "3alscKs" : $signed(forvar220))))};
              reg254 <= $unsigned(($signed(forvar238[(1'h0):(1'h0)]) <<< ("fR5" ?
                  reg184 : $signed($unsigned(reg236)))));
              reg255 = reg171;
              reg256 <= forvar238;
            end
        end
      else
        begin
          for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
            begin
              reg244 <= forvar209;
            end
          reg245 <= (((reg196[(4'h9):(2'h3)] && (-reg252)) * reg232[(4'hc):(3'h6)]) < "xFMiedQo5THpUMR");
        end
    end
  assign wire257 = $signed({$signed(($unsigned((8'hac)) ?
                           (reg171 << forvar178) : (wire136 || reg142)))});
  assign wire258 = {(forvar157[(1'h0):(1'h0)] && (8'hb0)),
                       (+{$unsigned(reg140), forvar203[(4'h9):(2'h3)]})};
  assign wire259 = reg222[(2'h3):(1'h0)];
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h8f9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire0;
  input wire signed [(5'h18):(1'h0)] wire1;
  input wire signed [(2'h3):(1'h0)] wire2;
  input wire [(4'hc):(1'h0)] wire3;
  input wire [(5'h13):(1'h0)] wire4;
  wire [(2'h2):(1'h0)] wire904;
  wire [(5'h16):(1'h0)] wire903;
  wire [(4'h8):(1'h0)] wire902;
  wire [(2'h3):(1'h0)] wire901;
  wire signed [(4'ha):(1'h0)] wire5;
  wire [(2'h2):(1'h0)] wire6;
  wire signed [(4'he):(1'h0)] wire60;
  wire [(5'h10):(1'h0)] wire61;
  wire [(5'h16):(1'h0)] wire79;
  wire signed [(5'h14):(1'h0)] wire843;
  wire signed [(4'h8):(1'h0)] wire845;
  wire [(4'hd):(1'h0)] wire846;
  wire signed [(4'hb):(1'h0)] wire857;
  wire [(4'he):(1'h0)] wire858;
  wire signed [(4'hd):(1'h0)] wire883;
  wire [(3'h6):(1'h0)] wire899;
  reg [(4'hb):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg9 = (1'h0);
  reg [(4'h8):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg13 = (1'h0);
  reg [(5'h18):(1'h0)] reg15 = (1'h0);
  reg [(3'h4):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg20 = (1'h0);
  reg [(2'h3):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg22 = (1'h0);
  reg [(4'hf):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg27 = (1'h0);
  reg [(5'h12):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg33 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg37 = (1'h0);
  reg [(4'hc):(1'h0)] reg39 = (1'h0);
  reg [(2'h2):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg41 = (1'h0);
  reg [(5'h12):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg43 = (1'h0);
  reg [(5'h15):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg52 = (1'h0);
  reg [(3'h4):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg57 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg62 = (1'h0);
  reg [(2'h2):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg69 = (1'h0);
  reg [(5'h17):(1'h0)] reg71 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg76 = (1'h0);
  reg signed [(4'he):(1'h0)] reg77 = (1'h0);
  reg [(5'h11):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg84 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg86 = (1'h0);
  reg [(5'h16):(1'h0)] reg88 = (1'h0);
  reg [(5'h18):(1'h0)] reg95 = (1'h0);
  reg [(5'h17):(1'h0)] reg97 = (1'h0);
  reg [(3'h4):(1'h0)] reg98 = (1'h0);
  reg [(4'h9):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg101 = (1'h0);
  reg [(4'ha):(1'h0)] reg103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg108 = (1'h0);
  reg [(4'h9):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg111 = (1'h0);
  reg [(3'h4):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg119 = (1'h0);
  reg [(2'h2):(1'h0)] reg848 = (1'h0);
  reg [(3'h4):(1'h0)] reg849 = (1'h0);
  reg [(5'h11):(1'h0)] reg850 = (1'h0);
  reg [(4'h8):(1'h0)] reg852 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg853 = (1'h0);
  reg [(5'h14):(1'h0)] reg854 = (1'h0);
  reg [(2'h2):(1'h0)] reg856 = (1'h0);
  reg [(3'h7):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg861 = (1'h0);
  reg [(5'h16):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg864 = (1'h0);
  reg [(3'h5):(1'h0)] reg871 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg873 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg876 = (1'h0);
  reg [(4'hb):(1'h0)] reg877 = (1'h0);
  reg [(5'h11):(1'h0)] reg881 = (1'h0);
  reg [(3'h4):(1'h0)] reg882 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg884 = (1'h0);
  reg [(5'h14):(1'h0)] reg885 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg886 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg895 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg897 = (1'h0);
  reg [(3'h7):(1'h0)] reg894 = (1'h0);
  reg [(5'h10):(1'h0)] reg893 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg892 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg891 = (1'h0);
  reg [(2'h3):(1'h0)] reg890 = (1'h0);
  reg [(3'h4):(1'h0)] forvar889 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg888 = (1'h0);
  reg [(4'hb):(1'h0)] forvar887 = (1'h0);
  reg [(3'h7):(1'h0)] reg880 = (1'h0);
  reg [(2'h2):(1'h0)] forvar879 = (1'h0);
  reg [(5'h17):(1'h0)] reg878 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar870 = (1'h0);
  reg [(3'h7):(1'h0)] forvar869 = (1'h0);
  reg [(5'h13):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg867 = (1'h0);
  reg [(3'h5):(1'h0)] forvar866 = (1'h0);
  reg [(3'h5):(1'h0)] reg865 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg863 = (1'h0);
  reg [(5'h17):(1'h0)] reg860 = (1'h0);
  reg [(5'h18):(1'h0)] reg855 = (1'h0);
  reg [(4'ha):(1'h0)] forvar847 = (1'h0);
  reg [(3'h7):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg847 = (1'h0);
  reg signed [(4'he):(1'h0)] reg118 = (1'h0);
  reg [(5'h14):(1'h0)] reg116 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar115 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar113 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar107 = (1'h0);
  reg [(5'h17):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg104 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg [(4'hb):(1'h0)] reg99 = (1'h0);
  reg [(5'h13):(1'h0)] reg96 = (1'h0);
  reg [(5'h10):(1'h0)] forvar94 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg92 = (1'h0);
  reg [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(5'h12):(1'h0)] reg90 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar89 = (1'h0);
  reg [(4'h8):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg85 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg81 = (1'h0);
  reg [(3'h7):(1'h0)] reg78 = (1'h0);
  reg [(5'h18):(1'h0)] reg75 = (1'h0);
  reg [(4'hb):(1'h0)] reg73 = (1'h0);
  reg [(4'hf):(1'h0)] reg70 = (1'h0);
  reg [(3'h7):(1'h0)] reg68 = (1'h0);
  reg [(4'h8):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg66 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg64 = (1'h0);
  reg [(4'hb):(1'h0)] reg63 = (1'h0);
  reg [(3'h6):(1'h0)] reg59 = (1'h0);
  reg [(5'h17):(1'h0)] forvar56 = (1'h0);
  reg [(2'h2):(1'h0)] reg55 = (1'h0);
  reg [(2'h2):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar49 = (1'h0);
  reg [(4'hd):(1'h0)] forvar48 = (1'h0);
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg38 = (1'h0);
  reg [(5'h18):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg35 = (1'h0);
  reg [(5'h10):(1'h0)] forvar34 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg30 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar29 = (1'h0);
  reg [(3'h7):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar15 = (1'h0);
  reg [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(5'h15):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar24 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar18 = (1'h0);
  reg [(5'h13):(1'h0)] forvar9 = (1'h0);
  reg [(4'hc):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg11 = (1'h0);
  assign y = {wire904,
                 wire903,
                 wire902,
                 wire901,
                 wire5,
                 wire6,
                 wire60,
                 wire61,
                 wire79,
                 wire843,
                 wire845,
                 wire846,
                 wire857,
                 wire858,
                 wire883,
                 wire899,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg12,
                 reg13,
                 reg15,
                 reg16,
                 reg17,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg27,
                 reg31,
                 reg33,
                 reg37,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 reg57,
                 reg58,
                 reg62,
                 reg65,
                 reg69,
                 reg71,
                 reg72,
                 reg74,
                 reg76,
                 reg77,
                 reg80,
                 reg83,
                 reg84,
                 reg86,
                 reg88,
                 reg95,
                 reg97,
                 reg98,
                 reg100,
                 reg101,
                 reg103,
                 reg105,
                 reg108,
                 reg109,
                 reg111,
                 reg112,
                 reg114,
                 reg117,
                 reg119,
                 reg848,
                 reg849,
                 reg850,
                 reg852,
                 reg853,
                 reg854,
                 reg856,
                 reg859,
                 reg861,
                 reg862,
                 reg864,
                 reg871,
                 reg872,
                 reg873,
                 reg876,
                 reg877,
                 reg881,
                 reg882,
                 reg884,
                 reg885,
                 reg886,
                 reg895,
                 reg896,
                 reg898,
                 reg897,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 forvar889,
                 reg888,
                 forvar887,
                 reg880,
                 forvar879,
                 reg878,
                 reg875,
                 reg874,
                 forvar870,
                 forvar869,
                 reg868,
                 reg867,
                 forvar866,
                 reg865,
                 reg863,
                 reg860,
                 reg855,
                 forvar847,
                 reg851,
                 reg847,
                 reg118,
                 reg116,
                 forvar115,
                 forvar113,
                 reg110,
                 forvar107,
                 reg106,
                 reg104,
                 reg102,
                 reg99,
                 reg96,
                 forvar94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 forvar89,
                 reg87,
                 reg85,
                 reg82,
                 reg81,
                 reg78,
                 reg75,
                 reg73,
                 reg70,
                 reg68,
                 reg67,
                 reg66,
                 reg64,
                 reg63,
                 reg59,
                 forvar56,
                 reg55,
                 reg54,
                 forvar49,
                 forvar48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg38,
                 reg36,
                 reg35,
                 forvar34,
                 reg32,
                 reg30,
                 forvar29,
                 reg18,
                 forvar15,
                 reg28,
                 reg26,
                 reg25,
                 forvar24,
                 reg19,
                 forvar18,
                 forvar9,
                 reg14,
                 reg11,
                 (1'h0)};
  assign wire5 = wire0[(4'hd):(3'h4)];
  assign wire6 = (wire1[(5'h16):(4'hf)] * wire0[(3'h4):(3'h4)]);
  always
    @(posedge clk) begin
      reg7 <= $unsigned(wire2);
      if ((wire0 ? (~^(~&$unsigned((^~wire1)))) : (8'hbc)))
        begin
          if ($unsigned({(wire4 >> ((^(8'h9e)) ? $unsigned(wire4) : wire0))}))
            begin
              reg8 <= $signed(wire1[(5'h17):(4'h9)]);
              reg9 <= (!((~&$unsigned(reg7)) ? (|wire4) : (8'ha2)));
              reg10 <= wire3;
              reg11 = {wire2[(1'h0):(1'h0)],
                  ({($signed(wire0) * {wire0})} ?
                      (^~wire3[(3'h5):(3'h4)]) : wire5[(3'h5):(3'h4)])};
              reg12 <= $signed(((reg8[(3'h6):(1'h0)] << (((8'hbb) - wire0) <= $unsigned(wire5))) + wire4));
            end
          else
            begin
              reg11 = $signed($unsigned(wire5));
              reg12 <= {reg11};
              reg13 <= reg10[(3'h5):(3'h4)];
              reg14 = ($signed($unsigned((-(+(8'ha6))))) >= reg7);
            end
        end
      else
        begin
          reg8 <= ((~^$signed(wire1)) << $signed((~$unsigned($signed(wire6)))));
          for (forvar9 = (1'h0); (forvar9 < (2'h3)); forvar9 = (forvar9 + (1'h1)))
            begin
              reg10 <= reg7[(1'h0):(1'h0)];
              reg12 <= ((!$signed($signed($signed(wire3)))) + $signed((~&$signed((~&wire0)))));
            end
        end
      if ((wire2 > reg11))
        begin
          reg15 <= $signed((^wire1[(5'h11):(4'ha)]));
          reg16 <= $unsigned($signed($signed($signed((^wire5)))));
          reg17 <= $signed(reg16);
          for (forvar18 = (1'h0); (forvar18 < (2'h3)); forvar18 = (forvar18 + (1'h1)))
            begin
              reg19 = reg17;
              reg20 <= $unsigned(({((8'ha9) ^~ reg7[(2'h2):(1'h1)]),
                  {(reg14 * wire4)}} || (+wire5)));
              reg21 <= (!forvar9[(5'h13):(3'h7)]);
              reg22 <= wire5;
              reg23 <= {((reg11[(3'h5):(1'h1)] | (^{wire2})) && reg19)};
            end
          for (forvar24 = (1'h0); (forvar24 < (1'h1)); forvar24 = (forvar24 + (1'h1)))
            begin
              reg25 = ($signed((-{$signed(reg9)})) ?
                  {$unsigned(reg13), reg19[(2'h3):(2'h2)]} : ((~({reg20, reg9} ?
                      (reg13 ?
                          (8'hbb) : reg14) : ((8'haa) == reg10))) ~^ {$unsigned($unsigned(reg22))}));
              reg26 = reg8[(3'h6):(3'h5)];
              reg27 <= $signed(reg17);
              reg28 = wire1[(5'h13):(1'h1)];
            end
        end
      else
        begin
          for (forvar15 = (1'h0); (forvar15 < (2'h3)); forvar15 = (forvar15 + (1'h1)))
            begin
              reg16 <= $signed($unsigned((~^(((8'h9c) ^~ reg13) ?
                  reg11[(5'h12):(5'h11)] : (reg21 ~^ reg27)))));
              reg18 = $unsigned(reg16[(1'h0):(1'h0)]);
              reg19 = reg9;
            end
          reg20 <= reg8[(4'ha):(4'h9)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar29 = (1'h0); (forvar29 < (1'h0)); forvar29 = (forvar29 + (1'h1)))
        begin
          if ((~&{reg23[(3'h7):(3'h6)]}))
            begin
              reg30 = reg27[(3'h7):(1'h0)];
            end
          else
            begin
              reg31 <= reg7;
              reg32 = $unsigned(reg8[(4'hb):(4'hb)]);
              reg33 <= reg15[(4'he):(4'h8)];
            end
        end
      for (forvar34 = (1'h0); (forvar34 < (2'h3)); forvar34 = (forvar34 + (1'h1)))
        begin
          reg35 = $unsigned(((reg32 && $signed($signed(wire1))) ?
              $unsigned($signed((reg10 < reg27))) : (reg16[(2'h2):(1'h1)] ?
                  (reg13 & (~&reg12)) : $signed(wire1))));
          if ((reg7[(1'h1):(1'h0)] ?
              (+$signed(($unsigned(wire4) ?
                  $unsigned(reg15) : (wire6 | wire4)))) : reg20))
            begin
              reg36 = ((-reg8[(2'h3):(2'h2)]) >= wire6[(1'h1):(1'h1)]);
            end
          else
            begin
              reg37 <= $signed($unsigned(($signed($unsigned(reg22)) * reg27)));
              reg38 = $signed((&$signed({$unsigned(reg31)})));
              reg39 <= {$unsigned($signed($signed(reg32))),
                  (({(|reg13), $unsigned(wire5)} ?
                          (wire5[(1'h0):(1'h0)] ?
                              reg13[(4'he):(4'hd)] : $signed(reg10)) : {$signed(reg33)}) ?
                      ((~(~(8'hb6))) ?
                          ({wire2, reg20} ?
                              (+reg31) : (reg32 ?
                                  forvar29 : reg38)) : $signed((&reg38))) : $unsigned((~$unsigned((8'hba)))))};
              reg40 <= ($signed({({reg17, reg31} <<< (reg27 ?
                      forvar34 : reg17))}) | $signed((~&(reg35[(3'h5):(1'h1)] ?
                  (~^wire4) : $unsigned(reg15)))));
            end
          if (reg17)
            begin
              reg41 <= ({(reg38 + ($signed((8'ha2)) < (~reg13)))} ?
                  $signed((reg22 ~^ $signed((~^reg15)))) : $signed($unsigned((~^$unsigned(reg7)))));
              reg42 <= {$signed(wire1),
                  $unsigned((((reg7 < reg17) <= (~(8'hb4))) ?
                      $unsigned(reg27[(4'hd):(4'h9)]) : $signed((!wire0))))};
              reg43 <= (~(!(({reg27} > wire0) | reg40)));
              reg44 = (reg36 <= reg13);
            end
          else
            begin
              reg41 <= wire4;
              reg42 <= reg27[(4'hd):(4'hc)];
              reg44 = (~&$signed(reg33[(3'h6):(1'h0)]));
              reg45 = $unsigned(reg32[(4'h8):(2'h2)]);
            end
          reg46 = (reg7 != (~^($signed(forvar29[(4'ha):(3'h6)]) || ({reg42,
                  wire2} ?
              (~reg45) : (reg37 ? wire1 : reg23)))));
          reg47 = $unsigned((7'h45));
        end
      for (forvar48 = (1'h0); (forvar48 < (2'h3)); forvar48 = (forvar48 + (1'h1)))
        begin
          for (forvar49 = (1'h0); (forvar49 < (2'h2)); forvar49 = (forvar49 + (1'h1)))
            begin
              reg50 <= $signed($unsigned(reg46[(4'hc):(1'h1)]));
            end
          if ($unsigned($unsigned(({(~^reg32),
              (reg23 ? reg50 : reg50)} >= forvar49[(2'h2):(1'h1)]))))
            begin
              reg51 <= ($signed($signed((reg44 ?
                      (wire1 != reg8) : ((8'ha9) ? reg7 : forvar49)))) ?
                  reg46 : {(-reg45),
                      (reg17[(1'h1):(1'h0)] ?
                          $signed({reg21}) : $unsigned((reg21 * wire1)))});
              reg52 <= {wire4[(4'hf):(2'h3)],
                  $unsigned(((forvar34 != $signed(forvar34)) && ({wire4} != (reg43 >>> reg39))))};
              reg53 <= reg40[(1'h0):(1'h0)];
            end
          else
            begin
              reg54 = $signed($unsigned($unsigned($signed($unsigned(reg52)))));
            end
          reg55 = (&($signed(reg51[(4'hc):(4'hc)]) ?
              $unsigned(reg13) : (~|$signed($unsigned(reg44)))));
          for (forvar56 = (1'h0); (forvar56 < (1'h1)); forvar56 = (forvar56 + (1'h1)))
            begin
              reg57 <= ($unsigned(reg31) ?
                  reg23 : $signed(((~forvar34) & ($unsigned(reg50) ?
                      $unsigned(reg17) : $signed(forvar49)))));
              reg58 <= reg20[(1'h1):(1'h0)];
            end
          reg59 = reg50[(5'h10):(4'he)];
        end
    end
  assign wire60 = reg7[(2'h3):(2'h2)];
  assign wire61 = reg20;
  always
    @(posedge clk) begin
      reg62 <= $unsigned((~|(reg17[(3'h4):(1'h0)] ? (!(reg9 | reg43)) : reg7)));
      if ((~reg42[(3'h7):(3'h4)]))
        begin
          reg63 = (((8'had) ? $unsigned(reg43) : {(~&(~&reg52))}) < reg27);
          if ($signed({{reg62, $unsigned((~|reg33))}}))
            begin
              reg64 = $unsigned((~|wire4));
              reg65 <= reg8[(4'ha):(2'h3)];
              reg66 = wire0[(2'h2):(1'h0)];
              reg67 = ($unsigned($signed($signed({reg23, reg10}))) ?
                  {(reg65 ? $signed((7'h42)) : reg8[(1'h0):(1'h0)]),
                      wire3[(3'h5):(2'h3)]} : ((~|(^~{(8'hb4),
                      wire0})) + {$unsigned(reg57[(2'h3):(2'h3)]),
                      (reg23 ?
                          (reg31 ? reg41 : reg58) : (reg57 ? reg22 : wire1))}));
            end
          else
            begin
              reg65 <= $signed((({(reg37 * reg16), reg13[(5'h13):(4'ha)]} ?
                  $signed(reg66[(3'h7):(3'h7)]) : (~&(reg66 << wire61))) < ({(~reg41)} ?
                  ((reg63 - wire3) > reg27[(4'hf):(4'hd)]) : ((~&(8'ha6)) ?
                      ((8'hbb) ^ reg57) : ((8'ha9) | (8'hbc))))));
            end
          if ($unsigned(reg58))
            begin
              reg68 = $unsigned($unsigned($signed((wire1[(4'h9):(1'h0)] ?
                  {reg50} : $unsigned(reg21)))));
            end
          else
            begin
              reg69 <= reg27;
              reg70 = $unsigned((^$signed($signed($unsigned(reg51)))));
            end
          if ($unsigned((reg42[(4'hf):(3'h7)] ?
              reg7[(2'h3):(2'h3)] : ($unsigned((reg51 > reg7)) >> (reg31 ?
                  reg8 : reg7[(3'h4):(2'h3)])))))
            begin
              reg71 <= {$signed(($unsigned(reg51) & reg33[(3'h6):(3'h6)]))};
              reg72 <= wire1[(3'h6):(2'h2)];
            end
          else
            begin
              reg71 <= (($unsigned({(wire61 ? reg31 : reg72)}) ?
                  (|($signed(reg43) ^~ (+reg70))) : wire61) >> (7'h41));
              reg72 <= (^$signed((-$unsigned(wire4[(1'h0):(1'h0)]))));
              reg73 = reg63;
              reg74 <= {reg71[(5'h14):(4'h8)]};
            end
          reg75 = {((({wire0, reg8} >>> (8'hb1)) * ((~|reg15) ?
                      {reg20, (7'h46)} : reg58)) ?
                  reg16[(1'h1):(1'h1)] : (~(~|((7'h44) ? reg52 : wire60)))),
              ((~|reg65) ?
                  $signed($unsigned($signed(wire0))) : $signed($signed($unsigned(reg10))))};
        end
      else
        begin
          if ({reg69[(4'h9):(2'h3)],
              (reg22[(3'h7):(3'h7)] ?
                  $signed($unsigned($signed(reg70))) : reg67[(3'h7):(3'h4)])})
            begin
              reg65 <= $signed($signed($unsigned({$signed(wire60),
                  $signed(wire5)})));
              reg69 <= $signed((~&(((!wire60) * $unsigned(reg57)) || reg52)));
              reg70 = reg15;
              reg73 = (-$unsigned((wire0[(4'hd):(3'h6)] ?
                  (~(^(8'ha1))) : ((^(8'hbd)) & $unsigned((8'h9f))))));
              reg75 = {reg42[(2'h3):(1'h0)]};
            end
          else
            begin
              reg65 <= (~(8'hb6));
              reg66 = $unsigned(reg74[(3'h4):(2'h2)]);
              reg69 <= (~&(($unsigned((~|reg72)) || reg52) ?
                  reg53[(2'h2):(2'h2)] : $signed(({wire61} & $signed(reg68)))));
              reg71 <= (($signed(reg23[(4'hd):(4'ha)]) ^~ $unsigned(reg42)) ?
                  reg8 : {$unsigned(((wire5 * (7'h49)) * (wire6 > reg63)))});
            end
          reg76 <= (~(~|{reg52}));
          reg77 <= reg31[(4'hd):(3'h5)];
          reg78 = (((reg40[(1'h1):(1'h0)] > ((reg33 ? reg76 : reg21) == (reg41 ?
                      wire3 : wire5))) ?
                  $signed($signed($unsigned(reg63))) : reg40) ?
              (|reg62) : (~&(^~reg63[(3'h7):(3'h4)])));
        end
    end
  assign wire79 = (!(reg33 || $unsigned({$signed(wire6), (wire0 && wire61)})));
  always
    @(posedge clk) begin
      reg80 <= {{reg69,
              $signed(($signed((8'hb1)) ? (reg7 <= (7'h42)) : (-reg69)))}};
      reg81 = (wire5[(3'h4):(2'h3)] ? reg62[(1'h1):(1'h0)] : reg16);
    end
  always
    @(posedge clk) begin
      if ((!$unsigned((~^$unsigned({reg7, wire4})))))
        begin
          reg82 = $signed($signed((reg76 ?
              ({(8'hab)} | ((7'h48) ? (8'hb6) : reg39)) : ((reg9 ?
                  wire60 : reg43) + (wire1 ? reg37 : (8'hb2))))));
        end
      else
        begin
          if ((+reg21))
            begin
              reg83 <= reg82;
              reg84 <= reg52[(5'h12):(4'h9)];
            end
          else
            begin
              reg82 = (|(+$unsigned({$unsigned(reg41)})));
              reg85 = ({(7'h42)} ^ $signed((!(reg58[(1'h1):(1'h1)] <<< {reg82}))));
              reg86 <= $unsigned(reg85);
              reg87 = reg43[(3'h5):(3'h4)];
              reg88 <= $unsigned((~&(reg12 - $signed((-wire4)))));
            end
          for (forvar89 = (1'h0); (forvar89 < (1'h1)); forvar89 = (forvar89 + (1'h1)))
            begin
              reg90 = (((~($unsigned(reg22) == (reg57 != reg7))) & $unsigned($unsigned((~&reg76)))) * (($signed($signed(reg80)) & reg8) >= $unsigned(($signed(reg10) ?
                  {reg43, (8'hb1)} : reg16))));
              reg91 = (~|reg40);
              reg92 = (((forvar89[(1'h1):(1'h1)] ?
                          forvar89 : wire4[(4'h9):(3'h7)]) ?
                      $unsigned((reg21[(2'h2):(1'h1)] ?
                          reg53 : $unsigned(reg82))) : $unsigned($unsigned($signed((8'hbe))))) ?
                  (reg20[(4'hf):(1'h0)] ?
                      (~^((wire60 ?
                          wire79 : wire61) + (reg8 <<< reg87))) : {(((7'h49) ?
                              reg77 : reg83) < $unsigned(reg88)),
                          $unsigned(wire79[(5'h15):(5'h10)])}) : reg84[(5'h10):(3'h6)]);
              reg93 = wire6[(1'h0):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar94 = (1'h0); (forvar94 < (2'h2)); forvar94 = (forvar94 + (1'h1)))
        begin
          if ((wire1 >= $unsigned((-$signed((|forvar94))))))
            begin
              reg95 <= reg22[(4'hd):(4'hc)];
              reg96 = {reg51};
            end
          else
            begin
              reg95 <= $signed(($signed($signed(reg7)) >= (^~wire5)));
              reg97 <= (^~$unsigned(wire6));
              reg98 <= $unsigned((reg9 ?
                  reg20 : ((8'h9e) ^ (&(wire3 ? reg51 : reg23)))));
            end
          reg99 = ((({reg16, (|reg72)} >>> $signed({(7'h46), reg12})) ?
              wire60 : $unsigned($unsigned(reg52))) ^~ reg72[(1'h1):(1'h1)]);
          if (reg9[(4'hf):(4'he)])
            begin
              reg100 <= (~|({(~|$signed(reg74)), (&$unsigned(reg39))} ?
                  wire2 : ($signed((reg37 ?
                      (7'h45) : wire3)) ^~ (~^reg21[(1'h1):(1'h1)]))));
              reg101 <= $unsigned((~&(reg16 + (^reg8))));
            end
          else
            begin
              reg100 <= ((8'hb0) ?
                  ((reg37 <<< ((reg88 || reg76) <<< $unsigned(wire1))) >>> (reg22[(1'h0):(1'h0)] ^~ reg12[(1'h1):(1'h0)])) : reg33);
              reg102 = (reg83[(3'h6):(1'h0)] ^~ $signed(reg100));
              reg103 <= (($signed((-{reg43})) ?
                      $signed($signed((reg62 ?
                          (8'hba) : reg41))) : (((^(8'hba)) ?
                          (^~reg15) : reg62) << (reg12[(2'h3):(2'h2)] > (reg86 == (7'h42))))) ?
                  (-(~|wire3)) : reg39);
              reg104 = {(((~^$unsigned(reg65)) >>> ({reg33, reg7} ?
                          (reg17 ? reg71 : wire1) : reg99[(2'h2):(1'h1)])) ?
                      (+((reg80 ? reg83 : wire79) ?
                          (^reg42) : (^reg103))) : ($unsigned($signed(reg74)) ?
                          $signed(reg37[(2'h3):(1'h1)]) : $signed($signed((8'hb4)))))};
            end
          reg105 <= ({$signed((reg76 ? {wire1} : $unsigned((8'hbb)))),
              ($signed((wire1 ?
                  reg17 : reg86)) * (+$unsigned(reg43)))} ^ reg33);
          reg106 = ({$unsigned({(reg52 ? reg37 : reg97),
                  (reg76 ? reg76 : reg88)}),
              ($signed(wire79) ?
                  $signed($signed(reg83)) : ($signed(wire2) ?
                      reg74[(4'h8):(2'h3)] : reg9))} + ($signed((&reg15[(5'h17):(3'h4)])) > $signed($signed((forvar94 + reg15)))));
        end
      for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
        begin
          reg108 <= $signed($unsigned($signed(((-reg106) ~^ reg102[(3'h6):(1'h1)]))));
          reg109 <= (+reg10);
          if ((!($signed(reg21) ? $unsigned(reg97) : (8'hbc))))
            begin
              reg110 = $signed((~^wire2));
              reg111 <= $unsigned($signed($unsigned((reg58[(3'h6):(1'h0)] | $unsigned((7'h48))))));
            end
          else
            begin
              reg110 = (~(reg20[(4'hc):(1'h1)] >> ($signed(wire4[(4'h8):(3'h6)]) ?
                  ($unsigned((7'h48)) ?
                      (reg96 || reg84) : (~(8'hb5))) : $unsigned(reg41[(5'h12):(3'h7)]))));
              reg111 <= (~|(^~$signed(((reg96 ^~ reg37) ?
                  reg40 : (reg57 - reg12)))));
              reg112 <= {(^$unsigned(reg40[(1'h1):(1'h1)]))};
            end
        end
      for (forvar113 = (1'h0); (forvar113 < (2'h3)); forvar113 = (forvar113 + (1'h1)))
        begin
          reg114 <= reg8;
          for (forvar115 = (1'h0); (forvar115 < (2'h3)); forvar115 = (forvar115 + (1'h1)))
            begin
              reg116 = reg80;
              reg117 <= (~&(8'h9c));
            end
          reg118 = {(reg20 ?
                  $signed((-(~wire6))) : $unsigned(forvar94[(2'h3):(1'h0)]))};
        end
      reg119 <= $signed($signed($unsigned((-$signed(reg16)))));
    end
  module120 #() modinst844 (.wire123(reg57), .wire122(reg8), .wire124(reg95), .y(wire843), .clk(clk), .wire121(reg76));
  assign wire845 = (+((((wire79 ? reg8 : reg22) ? $signed(reg9) : reg37) ?
                       (+$unsigned(reg52)) : (reg111[(4'ha):(3'h4)] < (wire60 ?
                           (8'ha1) : reg83))) == (!((reg77 & reg74) ?
                       $signed(reg7) : (^(8'ha4))))));
  assign wire846 = $signed(reg8[(5'h11):(1'h0)]);
  always
    @(posedge clk) begin
      if (((^{{((8'hbb) ? wire5 : (7'h48))},
          $unsigned($unsigned(reg71))}) && wire2))
        begin
          reg847 = reg88[(5'h13):(5'h10)];
          reg848 <= $unsigned($unsigned(reg16[(1'h0):(1'h0)]));
          if ($unsigned(($unsigned({reg58}) ?
              $unsigned(($signed(reg39) ?
                  $unsigned(reg50) : $signed(reg95))) : ((reg95 || reg8[(4'h8):(3'h7)]) != $signed($unsigned(reg57))))))
            begin
              reg849 <= ((reg74[(1'h1):(1'h1)] ?
                  $signed(($unsigned(reg16) ?
                      (~&reg41) : (&reg98))) : reg108[(4'h8):(2'h2)]) <<< {(+$signed($unsigned((7'h41))))});
              reg850 <= reg95[(5'h18):(5'h15)];
            end
          else
            begin
              reg849 <= {$unsigned({reg51, reg72[(2'h2):(2'h2)]})};
              reg850 <= wire846[(4'hd):(4'h8)];
            end
          reg851 = (($unsigned(reg10[(3'h4):(2'h2)]) ?
                  (reg12 ?
                      reg15[(5'h14):(4'he)] : $unsigned((reg111 ?
                          reg33 : wire6))) : (($signed(reg33) ?
                          wire3 : reg112[(3'h4):(2'h2)]) ?
                      $signed(wire61[(3'h5):(1'h0)]) : reg119[(1'h0):(1'h0)])) ?
              reg8 : (8'ha1));
        end
      else
        begin
          for (forvar847 = (1'h0); (forvar847 < (3'h4)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg851 = $signed(reg849[(3'h4):(1'h0)]);
            end
          reg852 <= ($unsigned(((reg8[(5'h11):(4'he)] << reg83[(5'h17):(2'h3)]) ?
                  {(reg71 ? reg40 : reg849)} : (~$signed(reg50)))) ?
              $unsigned(($unsigned((reg33 | reg112)) ?
                  $unsigned(reg8[(2'h3):(2'h3)]) : $signed($unsigned((8'hbc))))) : $signed((^~(~&(reg100 ?
                  reg105 : (8'h9c))))));
          reg853 <= $unsigned(((reg20[(5'h15):(3'h6)] < ({reg33, reg50} ?
              $signed(reg100) : wire5)) ~^ ((8'hb1) ?
              $unsigned((reg20 << reg40)) : ($signed(reg83) ?
                  (wire843 ^~ reg62) : {reg74}))));
          if ($unsigned(reg9[(4'hf):(4'h9)]))
            begin
              reg854 <= $unsigned($unsigned({((reg10 >= reg95) ?
                      wire845[(2'h3):(1'h1)] : reg848)}));
            end
          else
            begin
              reg855 = $unsigned($signed($signed($signed((reg83 ^~ (7'h44))))));
              reg856 <= reg42[(4'h8):(2'h2)];
            end
        end
    end
  assign wire857 = $signed(($unsigned({(~&reg16), reg88}) ?
                       reg83 : $signed($unsigned((reg848 ? reg50 : reg8)))));
  assign wire858 = reg37;
  always
    @(posedge clk) begin
      if ((~|((~|$signed((reg72 == (8'h9d)))) - (((wire4 ? reg100 : reg86) ?
              (|(8'ha5)) : $signed(reg62)) ?
          $unsigned((&reg50)) : (8'hb9)))))
        begin
          if ($unsigned((reg65 < $unsigned(reg74[(3'h7):(2'h2)]))))
            begin
              reg859 <= {(|reg7[(3'h5):(2'h3)]), reg42[(1'h0):(1'h0)]};
              reg860 = $signed($unsigned($signed(($signed(wire858) ~^ reg31))));
              reg861 <= ((reg40[(2'h2):(1'h0)] - $signed((|$unsigned(reg74)))) | (wire3[(4'hb):(1'h1)] ?
                  wire0[(2'h3):(2'h3)] : $signed(reg114[(1'h0):(1'h0)])));
              reg862 <= (^{(^~(reg22[(1'h0):(1'h0)] ^ reg850[(4'he):(4'hc)]))});
            end
          else
            begin
              reg860 = reg112[(2'h3):(2'h3)];
              reg863 = (!$signed(reg852[(4'h8):(3'h4)]));
            end
          reg864 <= reg42[(2'h2):(2'h2)];
        end
      else
        begin
          if (((^~reg861[(2'h2):(1'h0)]) ^ ((!$unsigned({reg862})) | $unsigned($unsigned(reg65)))))
            begin
              reg860 = $signed((-(reg33[(1'h1):(1'h1)] ?
                  ($unsigned((8'ha2)) ?
                      (~|(7'h49)) : (reg856 ? reg22 : reg860)) : (reg98 ?
                      (wire846 << reg850) : (!reg854)))));
              reg861 <= $signed((-reg849[(3'h4):(2'h2)]));
              reg862 <= $signed((reg41[(3'h4):(1'h1)] < (-(wire858[(4'h8):(2'h2)] ?
                  ((8'hb7) >= reg41) : reg9[(4'hc):(1'h0)]))));
            end
          else
            begin
              reg860 = (reg42[(5'h10):(5'h10)] ?
                  ((^~reg62) ?
                      wire846 : $unsigned(reg41[(3'h6):(1'h1)])) : reg76);
              reg861 <= $unsigned((-$signed(reg9[(4'h8):(1'h0)])));
              reg862 <= (wire845 <= reg52[(4'h9):(1'h0)]);
              reg864 <= reg72[(2'h3):(2'h2)];
            end
          reg865 = (~(~^$unsigned((-$signed(reg862)))));
          for (forvar866 = (1'h0); (forvar866 < (2'h2)); forvar866 = (forvar866 + (1'h1)))
            begin
              reg867 = $signed({(~(~&$signed((8'hae))))});
              reg868 = (reg65 != ((($signed(reg12) ?
                  (reg7 ? reg42 : (7'h42)) : (reg105 ?
                      reg97 : reg23)) <<< {((8'hb9) ?
                      reg860 : wire5)}) ~^ $unsigned((~$signed(reg10)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar869 = (1'h0); (forvar869 < (3'h4)); forvar869 = (forvar869 + (1'h1)))
        begin
          for (forvar870 = (1'h0); (forvar870 < (2'h2)); forvar870 = (forvar870 + (1'h1)))
            begin
              reg871 <= $signed($unsigned($unsigned(reg9)));
              reg872 <= reg101;
            end
          reg873 <= ((8'hb4) ?
              {(wire0[(1'h1):(1'h0)] >= {((8'hb6) ? reg103 : reg77)}),
                  $unsigned(($signed((8'ha5)) ~^ {reg40,
                      reg76}))} : reg8[(5'h10):(4'h8)]);
          if (($signed(((+$signed(reg27)) * (^~(reg69 >> reg86)))) ?
              {$unsigned(($unsigned(reg20) > wire61))} : (reg849[(3'h4):(2'h2)] ?
                  reg109 : (~^wire4[(5'h10):(4'hc)]))))
            begin
              reg874 = (reg105 ? (+(^~(|(~(8'hab))))) : reg77[(4'he):(3'h7)]);
              reg875 = $signed({{($signed(reg77) ?
                          (^~reg23) : reg111[(2'h2):(1'h0)])},
                  (((reg57 == (8'hb0)) == $unsigned(reg84)) ^~ $unsigned((reg112 ?
                      reg52 : reg7)))});
            end
          else
            begin
              reg874 = (($signed(wire843[(3'h4):(2'h2)]) && ($unsigned($unsigned(reg69)) << $unsigned(reg861))) ?
                  {$signed(((reg850 || reg84) >> (^~wire843))),
                      ($signed($signed(wire845)) ~^ reg864)} : ($signed(((^~wire857) ?
                          (!reg874) : (+wire0))) ?
                      $unsigned(reg80) : (~|$signed((-(8'h9d))))));
              reg876 <= $unsigned((&(8'hae)));
              reg877 <= $unsigned(($signed((~&(reg52 == reg43))) ?
                  (wire1 == ((^~forvar869) ?
                      (+reg111) : (~&reg27))) : reg856[(2'h2):(1'h0)]));
            end
          reg878 = (!$signed((reg21 ?
              wire79[(4'h9):(4'h9)] : (^~(reg86 ? forvar870 : reg13)))));
          for (forvar879 = (1'h0); (forvar879 < (2'h3)); forvar879 = (forvar879 + (1'h1)))
            begin
              reg880 = $signed((((|(reg859 ?
                  reg119 : (8'ha0))) <<< reg21) < forvar870[(3'h6):(3'h4)]));
              reg881 <= ($unsigned({(~(wire2 >>> wire4))}) ?
                  $signed(reg97[(4'hf):(4'ha)]) : reg62);
              reg882 <= (~&{((~^$signed((8'hb0))) && $unsigned($unsigned((8'had)))),
                  wire846[(3'h6):(1'h1)]});
            end
        end
    end
  assign wire883 = $signed((~&(reg37[(4'h8):(2'h3)] ?
                       reg111[(3'h5):(2'h2)] : $signed($signed(reg65)))));
  always
    @(posedge clk) begin
      reg884 <= reg861[(4'ha):(3'h6)];
      reg885 <= {((&{((8'ha9) | reg13), (wire3 ? reg848 : (8'had))}) ?
              $signed((((7'h40) ? reg872 : reg57) ?
                  $unsigned(reg856) : (reg10 ?
                      (8'ha0) : reg83))) : $unsigned({(reg862 ?
                      (8'h9d) : wire843),
                  (~|reg882)}))};
      reg886 <= ($signed((~reg119[(1'h1):(1'h1)])) ?
          (-$unsigned(reg39)) : reg57);
      for (forvar887 = (1'h0); (forvar887 < (1'h1)); forvar887 = (forvar887 + (1'h1)))
        begin
          reg888 = ($unsigned(reg41) ?
              $signed($signed($signed($unsigned(reg77)))) : wire883[(4'hb):(3'h5)]);
          for (forvar889 = (1'h0); (forvar889 < (2'h2)); forvar889 = (forvar889 + (1'h1)))
            begin
              reg890 = reg881[(4'hf):(4'hd)];
              reg891 = (wire4[(3'h6):(2'h3)] & reg21);
            end
          reg892 = reg37;
          reg893 = ({(($signed(reg9) * (~^reg848)) ~^ (reg119 <= reg111[(2'h2):(1'h0)]))} << (~&$unsigned((~|$signed(reg859)))));
          if ((((($signed((8'hb6)) + (^reg849)) ~^ {((7'h41) ^~ wire4)}) ?
              $signed(reg108[(3'h5):(3'h4)]) : (~&reg864[(5'h10):(2'h3)])) < $unsigned((+{(~(7'h47)),
              (wire858 ? reg12 : reg77)}))))
            begin
              reg894 = ({$signed(reg22)} >= ((((wire79 + (8'ha2)) ?
                      (reg108 ? (8'hb7) : reg856) : (reg58 - wire858)) ?
                  $signed($signed(reg861)) : (reg117[(3'h7):(1'h0)] ?
                      $unsigned(reg98) : (&wire60))) > reg114[(3'h5):(1'h0)]));
            end
          else
            begin
              reg895 <= $signed($signed(reg119));
              reg896 <= $unsigned($unsigned(reg95));
              reg897 = reg117;
              reg898 <= reg856[(1'h0):(1'h0)];
            end
        end
    end
  module125 #() modinst900 (.wire129(reg27), .y(wire899), .wire128(wire845), .wire127(reg42), .clk(clk), .wire126(reg88));
  assign wire901 = $unsigned($unsigned(((~&((7'h41) ^~ (8'hb8))) ?
                       (reg21[(2'h2):(1'h1)] ?
                           (reg849 * reg861) : reg62[(4'hb):(1'h0)]) : (7'h4a))));
  assign wire902 = $unsigned($unsigned(reg886));
  assign wire903 = wire901[(2'h2):(1'h1)];
  assign wire904 = (reg861 << reg877[(1'h1):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module120
#(parameter param842 = ((({{(8'ha2)}} ? {{(8'hac), (8'hb8)}, ((8'hb4) > (8'hb9))} : ((~(7'h48)) ? (-(7'h41)) : (~&(8'hae)))) ? (8'hbc) : ((^(~&(7'h47))) ? (((8'h9d) == (8'ha6)) << ((7'h47) ? (8'hb7) : (8'ha9))) : {{(8'ha7), (8'h9d)}, (8'hbd)})) ~^ (((^(8'hbc)) ? ((-(8'hba)) ? ((8'hb1) ? (8'hb2) : (8'ha4)) : ((8'h9e) ? (8'hb2) : (8'hb3))) : (((8'ha5) > (8'hba)) || ((8'hac) <= (8'h9c)))) ? (7'h40) : {(8'ha6)})))
(y, clk, wire124, wire123, wire122, wire121);
  output wire [(32'h3fa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire124;
  input wire signed [(4'hf):(1'h0)] wire123;
  input wire signed [(5'h17):(1'h0)] wire122;
  input wire [(4'he):(1'h0)] wire121;
  wire signed [(5'h11):(1'h0)] wire841;
  wire signed [(5'h17):(1'h0)] wire830;
  wire [(5'h12):(1'h0)] wire426;
  wire signed [(5'h12):(1'h0)] wire246;
  wire [(5'h15):(1'h0)] wire245;
  wire [(4'h9):(1'h0)] wire243;
  reg signed [(5'h16):(1'h0)] reg840 = (1'h0);
  reg [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg838 = (1'h0);
  reg [(5'h14):(1'h0)] reg837 = (1'h0);
  reg [(3'h7):(1'h0)] reg836 = (1'h0);
  reg [(4'hc):(1'h0)] reg835 = (1'h0);
  reg [(4'ha):(1'h0)] reg833 = (1'h0);
  reg [(2'h3):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg286 = (1'h0);
  reg [(5'h17):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg269 = (1'h0);
  reg [(3'h7):(1'h0)] reg267 = (1'h0);
  reg [(5'h10):(1'h0)] reg253 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg258 = (1'h0);
  reg [(4'h8):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg250 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg429 = (1'h0);
  reg [(4'hd):(1'h0)] reg430 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg [(5'h11):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg439 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg834 = (1'h0);
  reg [(5'h17):(1'h0)] forvar832 = (1'h0);
  reg [(4'ha):(1'h0)] reg438 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg436 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar435 = (1'h0);
  reg [(5'h16):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg428 = (1'h0);
  reg [(5'h14):(1'h0)] reg285 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar284 = (1'h0);
  reg [(3'h4):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg282 = (1'h0);
  reg [(5'h10):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar277 = (1'h0);
  reg [(5'h16):(1'h0)] reg276 = (1'h0);
  reg [(3'h7):(1'h0)] forvar275 = (1'h0);
  reg [(5'h17):(1'h0)] reg274 = (1'h0);
  reg [(3'h4):(1'h0)] reg271 = (1'h0);
  reg [(5'h17):(1'h0)] forvar270 = (1'h0);
  reg [(4'hc):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg266 = (1'h0);
  reg [(2'h2):(1'h0)] reg265 = (1'h0);
  reg [(4'hc):(1'h0)] forvar264 = (1'h0);
  reg [(5'h12):(1'h0)] reg263 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar262 = (1'h0);
  reg [(4'h9):(1'h0)] reg261 = (1'h0);
  reg [(4'hf):(1'h0)] reg260 = (1'h0);
  reg [(5'h14):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar257 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg256 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg254 = (1'h0);
  reg [(5'h18):(1'h0)] forvar253 = (1'h0);
  reg [(5'h10):(1'h0)] reg252 = (1'h0);
  reg signed [(4'he):(1'h0)] reg251 = (1'h0);
  reg [(3'h4):(1'h0)] forvar247 = (1'h0);
  assign y = {wire841,
                 wire830,
                 wire426,
                 wire246,
                 wire245,
                 wire243,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg833,
                 reg287,
                 reg286,
                 reg280,
                 reg279,
                 reg278,
                 reg273,
                 reg272,
                 reg269,
                 reg267,
                 reg253,
                 reg258,
                 reg257,
                 reg255,
                 reg250,
                 reg249,
                 reg248,
                 reg429,
                 reg430,
                 reg433,
                 reg434,
                 reg437,
                 reg439,
                 reg834,
                 forvar832,
                 reg438,
                 reg436,
                 forvar435,
                 reg432,
                 forvar431,
                 reg428,
                 reg285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 forvar277,
                 reg276,
                 forvar275,
                 reg274,
                 reg271,
                 forvar270,
                 reg268,
                 reg266,
                 reg265,
                 forvar264,
                 reg263,
                 forvar262,
                 reg261,
                 reg260,
                 reg259,
                 forvar257,
                 reg256,
                 reg254,
                 forvar253,
                 reg252,
                 reg251,
                 forvar247,
                 (1'h0)};
  module125 #() modinst244 (wire243, clk, wire121, wire123, wire124, wire122);
  assign wire245 = (7'h4a);
  assign wire246 = (^~(wire124[(3'h7):(2'h2)] == wire122));
  always
    @(posedge clk) begin
      if ((wire121 ?
          {wire124,
              (wire245[(4'he):(3'h5)] ?
                  $signed((wire121 ^ wire124)) : (wire122 ~^ {wire245,
                      (8'h9e)}))} : $signed(($unsigned(wire245[(4'hd):(3'h7)]) <= $unsigned((~|(8'hbd)))))))
        begin
          for (forvar247 = (1'h0); (forvar247 < (2'h2)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= ((^$signed(forvar247)) ? forvar247 : (~&wire123));
              reg249 <= $unsigned(({$signed((wire245 >> forvar247)),
                      forvar247[(3'h4):(2'h3)]} ?
                  {(wire123 ^ (wire243 ? wire124 : (8'hb1))),
                      ($unsigned(wire246) >>> $signed(wire122))} : wire123));
              reg250 <= $signed($unsigned(reg249[(3'h5):(3'h4)]));
              reg251 = ({(~|($unsigned(reg248) ?
                      (reg250 == wire122) : (reg249 << wire124)))} << (~(8'hbe)));
            end
          reg252 = (~&{$signed((wire245 ?
                  ((8'ha5) ? wire243 : reg248) : $signed(reg248)))});
          for (forvar253 = (1'h0); (forvar253 < (1'h0)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 = $signed((wire122[(2'h3):(2'h3)] ?
                  $unsigned(((wire124 > reg248) ?
                      reg249[(1'h0):(1'h0)] : $signed(reg248))) : $unsigned(wire243[(2'h3):(1'h1)])));
              reg255 <= wire245;
              reg256 = (~^wire246);
              reg257 <= (8'ha0);
              reg258 <= forvar253[(4'ha):(4'h8)];
            end
        end
      else
        begin
          for (forvar247 = (1'h0); (forvar247 < (2'h3)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= $unsigned(reg258[(2'h3):(2'h2)]);
              reg251 = (^~(~&$signed((-$signed(reg255)))));
              reg253 <= ($unsigned(wire122[(5'h11):(5'h11)]) > ({reg255,
                      wire245} ?
                  $signed(reg251) : wire123[(4'ha):(3'h4)]));
              reg255 <= (wire123 && (reg257[(2'h2):(2'h2)] ?
                  $signed(reg257) : ({$unsigned(reg254)} ?
                      $signed((reg258 ^ reg249)) : forvar253[(5'h13):(4'h9)])));
            end
          reg256 = (+wire243[(3'h7):(2'h3)]);
          for (forvar257 = (1'h0); (forvar257 < (2'h2)); forvar257 = (forvar257 + (1'h1)))
            begin
              reg259 = $unsigned(reg255);
              reg260 = reg248;
              reg261 = reg259;
            end
        end
      for (forvar262 = (1'h0); (forvar262 < (3'h4)); forvar262 = (forvar262 + (1'h1)))
        begin
          reg263 = (+reg256[(3'h7):(3'h4)]);
          for (forvar264 = (1'h0); (forvar264 < (1'h0)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 = $unsigned(reg254);
              reg266 = ($unsigned({(+$signed(reg248)),
                  ($signed(reg253) ~^ reg250[(4'hb):(1'h1)])}) + ((-reg249) ?
                  {(reg265 == {(8'hba), wire122}),
                      wire121[(4'he):(2'h2)]} : (^~(~&reg252))));
              reg267 <= reg252[(5'h10):(1'h0)];
              reg268 = (($unsigned((((8'hb5) ? wire124 : reg255) ^ ((8'h9f) ?
                      reg267 : wire243))) ^ (~(+wire124))) ?
                  reg261[(3'h5):(1'h1)] : forvar257);
              reg269 <= (forvar257 ?
                  {$unsigned($unsigned(reg267[(1'h1):(1'h1)]))} : (|((-reg261) ?
                      $unsigned(((8'h9f) && (7'h47))) : wire245)));
            end
          for (forvar270 = (1'h0); (forvar270 < (1'h1)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 = $unsigned(forvar253[(2'h2):(2'h2)]);
              reg272 <= ((reg250[(2'h2):(1'h0)] ?
                  (reg257[(2'h2):(1'h1)] | ($unsigned((8'ha6)) ?
                      (!reg258) : ((7'h44) ?
                          reg271 : wire246))) : $signed(forvar270)) == $unsigned($unsigned({$unsigned((8'ha3)),
                  forvar247})));
              reg273 <= ($signed($unsigned((-{wire123, reg266}))) ?
                  $signed(reg257) : ($unsigned((8'hb6)) ?
                      ($unsigned((reg256 ? (8'ha7) : reg254)) ?
                          $unsigned($signed(reg250)) : $unsigned(wire123)) : {$signed($signed(forvar270))}));
              reg274 = $signed(reg256[(5'h11):(4'h8)]);
            end
          for (forvar275 = (1'h0); (forvar275 < (2'h2)); forvar275 = (forvar275 + (1'h1)))
            begin
              reg276 = ($unsigned((~&((&forvar270) ?
                  (|reg258) : $unsigned(reg267)))) > wire123);
            end
        end
      for (forvar277 = (1'h0); (forvar277 < (3'h4)); forvar277 = (forvar277 + (1'h1)))
        begin
          reg278 <= (&(($signed($unsigned(reg261)) && reg258) ?
              (8'hb2) : $unsigned(((wire121 <= reg266) >>> reg273))));
          if (((-(-reg271[(2'h2):(1'h0)])) >= ($signed({wire124}) ?
              reg250 : $signed(($signed(forvar277) << (reg271 || forvar247))))))
            begin
              reg279 <= (~&wire121);
              reg280 <= (^~reg261);
              reg281 = $unsigned((reg251 ^ (7'h46)));
              reg282 = (^~$unsigned(reg259));
            end
          else
            begin
              reg279 <= $unsigned(((~&((+reg259) ? {reg250} : (~|reg267))) ?
                  $signed((+$signed((7'h43)))) : {$signed({(8'ha1)})}));
              reg281 = (reg254 ?
                  $signed((forvar253[(5'h18):(3'h5)] ?
                      $signed(reg282) : (^~(+reg260)))) : $unsigned(({(reg261 >> reg251),
                      $signed(forvar277)} == $unsigned($signed(wire124)))));
              reg282 = $signed(reg263[(4'ha):(2'h2)]);
              reg283 = $signed(($unsigned((~&$unsigned((8'hb4)))) ?
                  $unsigned($signed(forvar277[(1'h0):(1'h0)])) : {reg251[(2'h3):(2'h2)],
                      (~|wire124[(4'h9):(2'h3)])}));
            end
          for (forvar284 = (1'h0); (forvar284 < (3'h4)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 = ($signed(wire245[(4'hc):(4'h9)]) ?
                  reg272 : $unsigned((~^{(reg260 ^ (8'hba)),
                      (reg281 - (8'ha7))})));
              reg286 <= {$signed(reg258[(4'hd):(1'h0)]), reg255[(1'h1):(1'h1)]};
              reg287 <= forvar257;
            end
        end
    end
  module288 #() modinst427 (.wire291(reg286), .y(wire426), .clk(clk), .wire290(reg267), .wire289(reg253), .wire292(reg280), .wire293(reg257));
  always
    @(posedge clk) begin
      reg428 = {wire246[(4'he):(3'h7)]};
      reg429 <= reg272;
      reg430 <= (~|(~reg279));
      for (forvar431 = (1'h0); (forvar431 < (3'h4)); forvar431 = (forvar431 + (1'h1)))
        begin
          reg432 = (reg258 >>> (!$signed(($unsigned((8'h9d)) | (reg249 ?
              reg430 : reg286)))));
          reg433 <= $unsigned($unsigned(wire243));
          reg434 <= reg279;
          for (forvar435 = (1'h0); (forvar435 < (3'h4)); forvar435 = (forvar435 + (1'h1)))
            begin
              reg436 = ($unsigned(((reg258 ?
                  $signed(reg430) : (~|wire246)) >= $unsigned(((8'h9e) ?
                  reg253 : forvar435)))) >> $unsigned($signed((~|(reg429 != reg250)))));
              reg437 <= (8'haf);
              reg438 = (((8'hbe) & $signed(((wire121 ^ reg287) ^~ (reg267 ?
                      forvar431 : wire122)))) ?
                  ($signed($unsigned((wire122 ? (7'h49) : wire124))) ?
                      $signed(wire124) : ($unsigned($unsigned(wire243)) ?
                          ((reg437 == reg279) >>> (+reg279)) : ((~|reg280) <= reg269))) : $signed(reg428));
            end
          reg439 <= reg272;
        end
    end
  module440 #() modinst831 (wire830, clk, reg248, reg286, reg280, reg279, reg255);
  always
    @(posedge clk) begin
      for (forvar832 = (1'h0); (forvar832 < (2'h2)); forvar832 = (forvar832 + (1'h1)))
        begin
          if (($signed(($signed((-reg439)) ?
              ($unsigned(reg280) - (|reg255)) : wire121[(1'h1):(1'h0)])) ~^ {{$signed($unsigned(wire121)),
                  reg269[(4'ha):(3'h6)]}}))
            begin
              reg833 <= (($signed((reg287 == forvar832)) ?
                      (8'h9f) : {$signed(reg273[(2'h2):(1'h0)]),
                          ($signed(reg269) ?
                              wire245 : (reg280 ? reg248 : wire245))}) ?
                  (8'ha6) : {reg272[(3'h6):(3'h4)],
                      $unsigned($unsigned(wire426))});
              reg834 = reg249[(2'h2):(1'h1)];
            end
          else
            begin
              reg833 <= wire245[(3'h7):(3'h5)];
              reg834 = {($unsigned((reg833[(4'h8):(3'h7)] ^ wire426[(4'he):(2'h2)])) + (reg434 ^ ((^~reg279) | $signed(reg257))))};
              reg835 <= wire124[(2'h3):(1'h1)];
              reg836 <= wire830;
              reg837 <= (+({((reg279 ? wire246 : reg278) ?
                      ((8'had) | reg439) : (reg267 ?
                          reg833 : reg429))} >= $unsigned(((&reg273) ?
                  (reg248 ? wire426 : wire124) : reg834))));
            end
        end
      reg838 <= (wire830[(1'h1):(1'h0)] ?
          reg253 : ({($unsigned((7'h4a)) | $unsigned(reg430)),
              (reg434 ?
                  {(8'hbf), reg279} : $unsigned(reg287))} || $signed(wire246)));
      reg839 <= (&$unsigned((|$unsigned(wire246))));
      reg840 <= $signed(wire121);
    end
  assign wire841 = (~&$unsigned(reg250));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module440
#(parameter param828 = ((((~^((8'ha3) ? (8'ha0) : (7'h47))) * ((+(7'h41)) ? ((8'h9c) ? (8'hb3) : (8'hbd)) : (^~(7'h42)))) ? (8'ha3) : ((~^((8'ha2) | (7'h4a))) ^~ (((7'h49) ? (8'hbd) : (8'ha4)) ? ((8'h9c) <<< (8'ha4)) : {(8'h9f)}))) ? {{((8'ha4) ? ((7'h44) ~^ (8'hae)) : {(8'ha2)})}, {(((8'hb5) <<< (8'h9f)) << ((8'hb3) - (8'h9f)))}} : (((((8'h9e) ~^ (7'h47)) >>> (^~(8'hba))) ? ((+(8'ha0)) ? {(8'hbb)} : ((8'h9f) ? (8'hae) : (8'hbb))) : (8'hbd)) ? (({(8'hb3)} > (|(7'h44))) ? (^((8'hb9) ? (8'hb6) : (8'h9e))) : (((8'ha5) >> (8'hb9)) <= {(7'h45)})) : (!({(8'h9e), (7'h4a)} ? (~(7'h49)) : ((8'ha5) ? (7'h47) : (8'ha4)))))), 
parameter param829 = (+param828))
(y, clk, wire445, wire444, wire443, wire442, wire441);
  output wire [(32'hda):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire445;
  input wire [(5'h14):(1'h0)] wire444;
  input wire [(4'hf):(1'h0)] wire443;
  input wire signed [(5'h14):(1'h0)] wire442;
  input wire signed [(5'h16):(1'h0)] wire441;
  wire [(5'h12):(1'h0)] wire827;
  wire signed [(5'h10):(1'h0)] wire800;
  wire signed [(5'h10):(1'h0)] wire694;
  wire [(4'hb):(1'h0)] wire802;
  wire [(4'hb):(1'h0)] wire825;
  reg signed [(4'hf):(1'h0)] reg704 = (1'h0);
  reg [(3'h4):(1'h0)] reg700 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg699 = (1'h0);
  reg [(5'h18):(1'h0)] reg698 = (1'h0);
  reg [(2'h2):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg703 = (1'h0);
  reg [(5'h17):(1'h0)] reg702 = (1'h0);
  reg [(5'h18):(1'h0)] reg701 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar697 = (1'h0);
  assign y = {wire827,
                 wire800,
                 wire694,
                 wire802,
                 wire825,
                 reg704,
                 reg700,
                 reg699,
                 reg698,
                 reg696,
                 reg703,
                 reg702,
                 reg701,
                 forvar697,
                 (1'h0)};
  module446 #() modinst695 (wire694, clk, wire441, wire443, wire445, wire442);
  always
    @(posedge clk) begin
      reg696 <= (|(~^(($unsigned((8'hae)) ? wire444 : $signed(wire442)) ?
          wire442[(2'h3):(2'h3)] : $unsigned($signed(wire443)))));
      for (forvar697 = (1'h0); (forvar697 < (2'h2)); forvar697 = (forvar697 + (1'h1)))
        begin
          if ((((wire444[(3'h4):(2'h2)] ?
                  (!(wire442 ? (7'h47) : wire444)) : $unsigned((7'h4a))) ?
              reg696 : ((wire442 ?
                  $signed(wire444) : $signed((8'hb0))) <<< wire442)) ~^ wire444))
            begin
              reg698 <= $unsigned((~&(8'had)));
              reg699 <= $signed(forvar697);
              reg700 <= {(wire442[(1'h1):(1'h0)] ?
                      (8'ha7) : {($signed(reg699) ^ {wire441, wire443}),
                          reg699[(3'h7):(1'h1)]}),
                  $unsigned(wire443)};
              reg701 = reg696[(2'h2):(2'h2)];
              reg702 = $signed(((wire444 ?
                      $signed(((8'ha3) ?
                          reg696 : forvar697)) : ((|wire442) < forvar697[(1'h1):(1'h1)])) ?
                  $signed(((wire445 + (8'hba)) ?
                      wire694 : (wire694 ?
                          forvar697 : wire443))) : $signed({(wire441 || (8'hb8)),
                      $signed(wire441)})));
            end
          else
            begin
              reg698 <= ($unsigned($signed($unsigned(reg701[(5'h14):(1'h1)]))) ?
                  $unsigned($unsigned(reg700[(2'h3):(2'h3)])) : $signed(wire444[(4'hf):(3'h5)]));
              reg701 = $signed({reg700});
            end
          reg703 = ((({wire445[(4'hd):(3'h4)], reg699[(4'h9):(3'h6)]} ?
                  ({wire441, wire445} ?
                      $signed(wire445) : (8'h9c)) : reg699[(5'h13):(1'h0)]) ?
              ($unsigned($signed(wire442)) >= $unsigned(forvar697)) : $unsigned({$signed(reg698),
                  (reg699 == wire444)})) || wire694[(3'h7):(2'h3)]);
        end
      reg704 <= ($signed({((wire443 ? reg703 : reg700) ?
                  $signed(wire441) : (^~wire444)),
              (((8'hbd) ? (8'hb1) : wire694) - (reg696 ~^ wire442))}) ?
          wire694[(4'hb):(1'h1)] : $unsigned((+({reg702} - {(8'hb8),
              wire445}))));
    end
  module705 #() modinst801 (.wire708(wire694), .clk(clk), .wire709(wire445), .y(wire800), .wire707(reg698), .wire706(wire442));
  assign wire802 = wire441[(5'h15):(1'h1)];
  module803 #() modinst826 (wire825, clk, wire442, wire800, reg699, wire694);
  assign wire827 = $unsigned(wire802);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module288  (y, clk, wire293, wire292, wire291, wire290, wire289);
  output wire [(32'h6c3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire293;
  input wire signed [(3'h5):(1'h0)] wire292;
  input wire signed [(2'h2):(1'h0)] wire291;
  input wire [(3'h7):(1'h0)] wire290;
  input wire [(4'ha):(1'h0)] wire289;
  wire signed [(5'h15):(1'h0)] wire424;
  wire signed [(5'h16):(1'h0)] wire420;
  wire [(2'h2):(1'h0)] wire361;
  wire signed [(4'he):(1'h0)] wire360;
  wire signed [(5'h10):(1'h0)] wire324;
  wire [(4'h8):(1'h0)] wire297;
  wire signed [(4'h9):(1'h0)] wire296;
  wire signed [(4'hb):(1'h0)] wire295;
  wire signed [(3'h5):(1'h0)] wire294;
  reg [(4'hf):(1'h0)] reg418 = (1'h0);
  reg [(4'he):(1'h0)] reg415 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg407 = (1'h0);
  reg [(5'h11):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg402 = (1'h0);
  reg [(5'h12):(1'h0)] reg396 = (1'h0);
  reg signed [(4'he):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg392 = (1'h0);
  reg [(2'h3):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg387 = (1'h0);
  reg [(3'h4):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg375 = (1'h0);
  reg [(3'h4):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg368 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg365 = (1'h0);
  reg [(5'h11):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg354 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg353 = (1'h0);
  reg [(5'h16):(1'h0)] reg347 = (1'h0);
  reg [(2'h3):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg346 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg344 = (1'h0);
  reg [(4'h8):(1'h0)] reg343 = (1'h0);
  reg [(4'hf):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg337 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg335 = (1'h0);
  reg [(5'h15):(1'h0)] reg332 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg331 = (1'h0);
  reg [(4'h9):(1'h0)] reg328 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg323 = (1'h0);
  reg [(3'h4):(1'h0)] reg321 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg318 = (1'h0);
  reg [(5'h15):(1'h0)] reg317 = (1'h0);
  reg [(5'h12):(1'h0)] reg314 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg312 = (1'h0);
  reg [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg306 = (1'h0);
  reg [(2'h3):(1'h0)] reg303 = (1'h0);
  reg [(3'h6):(1'h0)] reg302 = (1'h0);
  reg [(5'h18):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg425 = (1'h0);
  reg [(5'h17):(1'h0)] reg423 = (1'h0);
  reg [(5'h13):(1'h0)] reg422 = (1'h0);
  reg [(4'h8):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg419 = (1'h0);
  reg [(3'h4):(1'h0)] reg417 = (1'h0);
  reg [(4'hb):(1'h0)] reg416 = (1'h0);
  reg [(4'h8):(1'h0)] reg413 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg411 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg410 = (1'h0);
  reg [(2'h2):(1'h0)] forvar409 = (1'h0);
  reg [(4'hb):(1'h0)] reg406 = (1'h0);
  reg [(4'hd):(1'h0)] reg405 = (1'h0);
  reg [(5'h18):(1'h0)] reg401 = (1'h0);
  reg [(5'h17):(1'h0)] reg400 = (1'h0);
  reg [(5'h14):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg397 = (1'h0);
  reg [(3'h4):(1'h0)] forvar395 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar394 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar389 = (1'h0);
  reg [(5'h11):(1'h0)] forvar388 = (1'h0);
  reg [(5'h15):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg385 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg384 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg383 = (1'h0);
  reg [(4'hf):(1'h0)] reg382 = (1'h0);
  reg [(4'hb):(1'h0)] reg381 = (1'h0);
  reg [(5'h11):(1'h0)] forvar380 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg378 = (1'h0);
  reg [(5'h12):(1'h0)] reg376 = (1'h0);
  reg [(5'h18):(1'h0)] forvar374 = (1'h0);
  reg [(2'h2):(1'h0)] reg373 = (1'h0);
  reg [(3'h6):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg371 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar369 = (1'h0);
  reg [(2'h2):(1'h0)] reg367 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg366 = (1'h0);
  reg [(5'h16):(1'h0)] forvar364 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg359 = (1'h0);
  reg [(2'h2):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg356 = (1'h0);
  reg [(2'h2):(1'h0)] reg352 = (1'h0);
  reg [(5'h12):(1'h0)] forvar351 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg348 = (1'h0);
  reg [(4'h8):(1'h0)] forvar347 = (1'h0);
  reg [(3'h6):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar340 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg336 = (1'h0);
  reg [(5'h17):(1'h0)] reg334 = (1'h0);
  reg [(4'ha):(1'h0)] forvar333 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg330 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg [(5'h11):(1'h0)] forvar327 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar326 = (1'h0);
  reg [(4'he):(1'h0)] reg325 = (1'h0);
  reg [(4'h8):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar316 = (1'h0);
  reg [(4'hf):(1'h0)] reg315 = (1'h0);
  reg [(4'h8):(1'h0)] reg313 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg311 = (1'h0);
  reg [(4'hf):(1'h0)] reg310 = (1'h0);
  reg signed [(4'he):(1'h0)] reg308 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar305 = (1'h0);
  reg [(5'h17):(1'h0)] forvar304 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar299 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg298 = (1'h0);
  assign y = {wire424,
                 wire420,
                 wire361,
                 wire360,
                 wire324,
                 wire297,
                 wire296,
                 wire295,
                 wire294,
                 reg418,
                 reg415,
                 reg414,
                 reg408,
                 reg407,
                 reg404,
                 reg403,
                 reg402,
                 reg396,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg387,
                 reg379,
                 reg377,
                 reg375,
                 reg372,
                 reg368,
                 reg365,
                 reg363,
                 reg362,
                 reg358,
                 reg355,
                 reg354,
                 reg353,
                 reg347,
                 reg350,
                 reg346,
                 reg344,
                 reg343,
                 reg339,
                 reg338,
                 reg337,
                 reg335,
                 reg332,
                 reg331,
                 reg328,
                 reg323,
                 reg321,
                 reg320,
                 reg318,
                 reg317,
                 reg314,
                 reg312,
                 reg309,
                 reg307,
                 reg306,
                 reg303,
                 reg302,
                 reg300,
                 reg425,
                 reg423,
                 reg422,
                 reg421,
                 reg419,
                 reg417,
                 reg416,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 forvar409,
                 reg406,
                 reg405,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 forvar395,
                 forvar394,
                 forvar389,
                 forvar388,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 forvar380,
                 reg378,
                 reg376,
                 forvar374,
                 reg373,
                 reg364,
                 reg371,
                 reg370,
                 forvar369,
                 reg367,
                 reg366,
                 forvar364,
                 reg359,
                 reg357,
                 reg356,
                 reg352,
                 forvar351,
                 reg349,
                 reg348,
                 forvar347,
                 reg345,
                 reg342,
                 reg341,
                 forvar340,
                 reg336,
                 reg334,
                 forvar333,
                 reg330,
                 reg329,
                 forvar327,
                 forvar326,
                 reg325,
                 reg322,
                 reg319,
                 forvar316,
                 reg315,
                 reg313,
                 reg311,
                 reg310,
                 reg308,
                 forvar305,
                 forvar304,
                 reg301,
                 forvar299,
                 reg298,
                 (1'h0)};
  assign wire294 = (~|wire289[(3'h6):(2'h2)]);
  assign wire295 = $signed({(({wire290, wire291} ?
                           (7'h40) : wire290) * {wire293[(1'h0):(1'h0)]})});
  assign wire296 = wire293;
  assign wire297 = (^~wire292[(3'h5):(2'h3)]);
  always
    @(posedge clk) begin
      reg298 = wire296;
      for (forvar299 = (1'h0); (forvar299 < (3'h4)); forvar299 = (forvar299 + (1'h1)))
        begin
          if (wire294)
            begin
              reg300 <= $unsigned(forvar299);
            end
          else
            begin
              reg301 = {wire294[(2'h3):(2'h3)]};
              reg302 <= (|(($signed(wire293[(2'h2):(2'h2)]) > $signed(wire297[(2'h3):(1'h1)])) ^~ (($signed((8'ha5)) >= (wire293 ?
                  (8'hb7) : (8'hb8))) & $signed(((8'hb0) < wire290)))));
            end
          reg303 <= $unsigned((reg302 ?
              $signed(((reg298 ? reg300 : wire289) ?
                  (-wire296) : {wire296})) : ($unsigned((~^wire291)) ?
                  wire291[(1'h0):(1'h0)] : ((reg298 ? wire292 : wire291) ?
                      (^~(8'hb3)) : reg301[(1'h1):(1'h0)]))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
        begin
          for (forvar305 = (1'h0); (forvar305 < (1'h1)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 <= (-(^~wire291));
              reg307 <= {$unsigned(((^wire295) ?
                      (^wire293) : forvar304[(2'h3):(2'h2)]))};
              reg308 = ({$unsigned((~reg306[(4'hb):(4'ha)]))} >> wire297);
              reg309 <= {$unsigned((-reg303[(1'h1):(1'h1)]))};
            end
          if ({{{$unsigned($signed(wire290)),
                      ((wire290 ? reg306 : forvar305) ?
                          (reg303 ^~ reg309) : (~&wire292))},
                  forvar304}})
            begin
              reg310 = {$signed(reg308)};
              reg311 = wire295;
              reg312 <= $signed(($unsigned(reg302[(3'h5):(3'h4)]) ~^ ($unsigned((wire290 <<< (7'h47))) ?
                  wire289[(3'h4):(3'h4)] : reg300)));
              reg313 = ((reg311[(1'h1):(1'h1)] | ($unsigned((8'hb9)) ?
                  {(wire296 ? wire294 : reg302), reg306} : ($unsigned(reg303) ?
                      reg307[(3'h6):(1'h0)] : $unsigned(wire296)))) * forvar304[(5'h17):(4'hc)]);
              reg314 <= $signed(reg309[(3'h4):(1'h1)]);
            end
          else
            begin
              reg310 = ((+(($unsigned(wire295) ?
                  (^~wire291) : wire295) == reg314[(2'h3):(1'h0)])) & reg309);
              reg312 <= $signed({reg314[(2'h3):(1'h0)], (~(&(+reg310)))});
              reg313 = $unsigned(((({wire289, (8'ha5)} ?
                      reg311 : wire296[(1'h0):(1'h0)]) && (^~$signed((7'h40)))) ?
                  ($unsigned(((8'ha5) ? wire290 : (8'hb6))) ?
                      $unsigned($signed(reg307)) : ((8'hbf) ?
                          (reg309 ?
                              wire290 : reg312) : reg314)) : (&reg307[(4'h8):(3'h4)])));
              reg315 = wire293;
            end
          for (forvar316 = (1'h0); (forvar316 < (1'h1)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 <= ($signed($signed(($unsigned(wire291) ^~ forvar305[(2'h3):(2'h3)]))) ?
                  $signed(($unsigned((forvar316 ? reg303 : reg314)) ?
                      reg314 : $unsigned((wire294 ?
                          (8'ha1) : (8'hb9))))) : (($signed((forvar305 ?
                              reg302 : reg308)) ?
                          $unsigned(reg310) : (!(wire290 | wire296))) ?
                      wire296[(1'h1):(1'h0)] : (reg313[(3'h7):(1'h1)] ?
                          (8'ha8) : ($unsigned(reg300) ?
                              (reg302 || wire297) : {reg313, reg312}))));
              reg318 <= $signed($signed(wire289[(4'h9):(2'h3)]));
              reg319 = ($signed($unsigned(reg306[(4'h8):(3'h7)])) ?
                  reg308[(4'h8):(1'h0)] : $signed({wire296}));
              reg320 <= $signed((~&(7'h40)));
              reg321 <= $unsigned(reg312[(3'h7):(2'h2)]);
            end
          reg322 = (reg313 ?
              ((8'hb4) ?
                  ($unsigned($signed(reg315)) >= (~{(8'hb8)})) : $signed(reg302[(2'h3):(2'h3)])) : $signed((reg318 >>> ($unsigned(reg307) ?
                  $unsigned(reg306) : ((8'hab) < reg317)))));
        end
      reg323 <= (&reg306);
    end
  assign wire324 = reg312[(2'h3):(2'h3)];
  always
    @(posedge clk) begin
      reg325 = $signed($unsigned(((^~reg312) ?
          $signed(reg314) : (^~$signed(reg312)))));
      for (forvar326 = (1'h0); (forvar326 < (3'h4)); forvar326 = (forvar326 + (1'h1)))
        begin
          for (forvar327 = (1'h0); (forvar327 < (3'h4)); forvar327 = (forvar327 + (1'h1)))
            begin
              reg328 <= wire292[(2'h2):(1'h0)];
              reg329 = (wire291[(1'h0):(1'h0)] >>> (~^reg306[(4'h8):(3'h4)]));
              reg330 = reg328;
              reg331 <= forvar326;
              reg332 <= (reg320 ? (~&(!$signed((-reg302)))) : wire290);
            end
          for (forvar333 = (1'h0); (forvar333 < (2'h3)); forvar333 = (forvar333 + (1'h1)))
            begin
              reg334 = (((wire290[(2'h3):(2'h3)] >= reg309) * $unsigned($signed((reg330 ?
                  reg318 : (8'h9e))))) < $signed(reg317));
              reg335 <= reg323;
              reg336 = (^$unsigned(wire290));
              reg337 <= $unsigned($signed(reg303[(1'h0):(1'h0)]));
            end
          reg338 <= reg306;
          reg339 <= reg309[(2'h3):(2'h2)];
          for (forvar340 = (1'h0); (forvar340 < (2'h3)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 = (((($signed(reg321) ?
                      {forvar340} : (wire324 ?
                          (8'hbc) : wire324)) + wire290[(3'h5):(2'h2)]) ?
                  (reg323 * ((&forvar326) ? reg332 : (+(8'hbf)))) : ((7'h41) ?
                      (&$signed(wire291)) : reg320[(3'h4):(1'h1)])) >> $unsigned(wire295));
              reg342 = (reg339[(3'h6):(3'h4)] ^~ $unsigned(wire292[(3'h5):(1'h1)]));
              reg343 <= ($unsigned(reg320[(3'h6):(3'h4)]) >> {{$signed((-wire297)),
                      (forvar340 ? $unsigned(reg309) : $unsigned((7'h43)))},
                  wire290});
              reg344 <= $signed(({$unsigned($unsigned(wire291)),
                      (reg331 != wire294)} ?
                  ({reg312[(1'h0):(1'h0)]} >> {reg338,
                      (reg342 ?
                          reg320 : reg342)}) : ((reg317[(4'hc):(3'h5)] < $signed((8'ha3))) + $signed((8'hae)))));
            end
        end
      reg345 = $unsigned(reg312);
      reg346 <= (reg314[(3'h5):(2'h3)] ?
          (wire289[(2'h3):(2'h3)] + ({(reg345 ? reg332 : wire324),
              $unsigned((7'h49))} > forvar340[(2'h3):(2'h2)])) : {({reg325,
                  reg336[(2'h3):(2'h3)]} >= {reg341,
                  (forvar333 ? reg300 : reg318)}),
              $unsigned(($signed((8'hb9)) ?
                  (reg344 ? reg306 : (7'h46)) : (reg343 > reg342)))});
      if (forvar327)
        begin
          for (forvar347 = (1'h0); (forvar347 < (2'h2)); forvar347 = (forvar347 + (1'h1)))
            begin
              reg348 = reg329[(2'h3):(2'h3)];
              reg349 = (({reg338, $unsigned((reg300 ? wire289 : reg341))} ?
                      (8'hab) : ((8'ha3) ^ (forvar340 + (reg318 <<< reg321)))) ?
                  $unsigned({$unsigned((reg346 ?
                          reg307 : reg300))}) : reg317[(4'hc):(2'h2)]);
              reg350 <= reg318;
            end
        end
      else
        begin
          if (reg346[(1'h1):(1'h1)])
            begin
              reg347 <= $signed((|(~^(~^$unsigned((8'ha3))))));
            end
          else
            begin
              reg347 <= $unsigned(((8'hbd) ? reg323 : $unsigned(reg341)));
              reg348 = wire324[(3'h6):(1'h1)];
              reg349 = $unsigned($unsigned({{(~|wire294)}}));
              reg350 <= ($unsigned(((+reg332) ?
                      {{reg312, reg344}} : (&(reg325 << (7'h40))))) ?
                  {reg334[(5'h17):(5'h17)], reg321} : reg331[(1'h0):(1'h0)]);
            end
          for (forvar351 = (1'h0); (forvar351 < (2'h3)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 = reg342[(5'h13):(4'ha)];
              reg353 <= (!(^$signed(reg344)));
              reg354 <= (~^(((((7'h46) >> (7'h41)) ? reg347 : (~&reg306)) ?
                  reg332 : ((8'hae) <<< (~&reg309))) >= reg347));
              reg355 <= $unsigned(reg328[(4'h8):(3'h5)]);
              reg356 = forvar347;
            end
          reg357 = ({(reg329 ?
                      ((^~reg325) >= (reg342 ?
                          wire293 : forvar351)) : (!(!forvar333))),
                  reg355[(2'h3):(1'h1)]} ?
              $signed({reg348, reg338}) : reg356);
          reg358 <= (-reg345);
        end
    end
  always
    @(posedge clk) begin
      reg359 = $unsigned(($signed(reg321) ~^ $signed($unsigned(reg338[(4'hd):(4'h8)]))));
    end
  assign wire360 = reg331[(3'h7):(1'h0)];
  assign wire361 = reg339;
  always
    @(posedge clk) begin
      if ({reg321,
          {($unsigned((^~reg355)) ?
                  reg358 : ($signed(reg312) ? (-reg335) : $signed(reg339))),
              $unsigned($unsigned((|(8'ha2))))}})
        begin
          reg362 <= reg347;
          reg363 <= wire324;
          for (forvar364 = (1'h0); (forvar364 < (1'h1)); forvar364 = (forvar364 + (1'h1)))
            begin
              reg365 <= $unsigned((~&wire292[(1'h0):(1'h0)]));
              reg366 = $unsigned($signed(reg303[(1'h1):(1'h0)]));
              reg367 = reg347;
            end
          reg368 <= reg320[(3'h5):(2'h3)];
          for (forvar369 = (1'h0); (forvar369 < (1'h0)); forvar369 = (forvar369 + (1'h1)))
            begin
              reg370 = ({reg344[(1'h1):(1'h0)]} > wire324[(4'hc):(3'h4)]);
              reg371 = reg332[(2'h3):(2'h2)];
              reg372 <= reg321;
            end
        end
      else
        begin
          reg362 <= $unsigned((&$unsigned(((^reg335) + $signed(wire295)))));
          reg363 <= reg371[(5'h10):(4'hb)];
          if ((({((reg335 ? reg358 : wire289) ?
                          ((7'h42) ? reg321 : reg346) : (wire324 >= reg347))} ?
                  reg347 : {reg314, reg306}) ?
              reg372 : $unsigned((+{(reg323 >> reg365),
                  wire291[(1'h1):(1'h0)]}))))
            begin
              reg364 = ($signed($unsigned(reg303[(2'h2):(1'h0)])) | wire292);
              reg366 = (((!($signed((8'hac)) < ((7'h48) <= reg358))) || reg337) || (|wire324));
            end
          else
            begin
              reg364 = reg318[(2'h2):(2'h2)];
              reg365 <= wire291;
              reg366 = $signed({((-reg371[(3'h7):(2'h2)]) || (reg303[(2'h2):(1'h1)] ?
                      $unsigned(reg343) : reg355[(3'h5):(1'h1)])),
                  ((~(8'hb9)) ? {(wire290 || reg354)} : reg363)});
            end
        end
      reg373 = {$unsigned($signed({{reg364}, (reg328 + reg307)})),
          ($signed(((+reg302) || reg365)) * $signed((+reg365)))};
      for (forvar374 = (1'h0); (forvar374 < (3'h4)); forvar374 = (forvar374 + (1'h1)))
        begin
          if ($unsigned(($signed($unsigned(reg306[(4'hc):(2'h3)])) != reg323)))
            begin
              reg375 <= wire360[(2'h3):(2'h2)];
              reg376 = reg320[(3'h4):(3'h4)];
              reg377 <= $unsigned((|$signed((reg337[(1'h1):(1'h0)] ?
                  $signed(reg375) : wire293[(1'h1):(1'h0)]))));
              reg378 = reg376[(1'h1):(1'h1)];
              reg379 <= reg364;
            end
          else
            begin
              reg375 <= reg353[(3'h5):(2'h2)];
              reg377 <= $signed($signed($unsigned($signed((^wire289)))));
              reg378 = (8'hb9);
            end
          for (forvar380 = (1'h0); (forvar380 < (2'h2)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 = $signed({$unsigned((|(wire297 ^ reg353)))});
              reg382 = (8'hb5);
              reg383 = {reg368};
              reg384 = reg376[(4'he):(3'h5)];
            end
        end
      reg385 = reg355[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg386 = reg335;
      reg387 <= $unsigned((+$unsigned(({reg320} != $unsigned(reg363)))));
      for (forvar388 = (1'h0); (forvar388 < (2'h2)); forvar388 = (forvar388 + (1'h1)))
        begin
          for (forvar389 = (1'h0); (forvar389 < (1'h0)); forvar389 = (forvar389 + (1'h1)))
            begin
              reg390 <= (&($signed($unsigned(reg355)) ?
                  reg363[(4'h8):(2'h3)] : {(|reg303[(1'h1):(1'h0)]),
                      (~&$signed(reg350))}));
              reg391 <= (&$unsigned(reg387));
              reg392 <= {($unsigned($unsigned($unsigned(reg347))) ?
                      $unsigned($unsigned({reg343,
                          reg307})) : $unsigned($signed(wire360[(3'h7):(2'h2)]))),
                  (~^(((reg300 ? reg332 : (8'ha0)) < $signed((8'hab))) ?
                      (~^reg379[(2'h2):(1'h1)]) : $unsigned((~&reg314))))};
              reg393 <= (~|wire293[(1'h1):(1'h0)]);
            end
        end
      for (forvar394 = (1'h0); (forvar394 < (2'h3)); forvar394 = (forvar394 + (1'h1)))
        begin
          for (forvar395 = (1'h0); (forvar395 < (3'h4)); forvar395 = (forvar395 + (1'h1)))
            begin
              reg396 <= $signed((8'ha1));
              reg397 = (reg328[(3'h6):(3'h5)] ~^ (~&(~$signed((~reg347)))));
              reg398 = wire291;
              reg399 = ({reg353[(1'h0):(1'h0)],
                      (reg362[(5'h13):(1'h1)] ?
                          $signed(reg377) : $signed(((8'ha5) || reg309)))} ?
                  reg306[(3'h6):(3'h4)] : reg320[(3'h4):(1'h1)]);
              reg400 = ((7'h43) ?
                  $signed(reg320[(2'h3):(2'h2)]) : $signed(forvar394[(3'h4):(1'h1)]));
            end
        end
      if (($unsigned(($signed((reg398 > reg320)) ?
          $unsigned((^reg368)) : (~(wire324 != reg302)))) || (($signed((~^reg398)) && (^~(reg377 - (8'h9c)))) ?
          (((reg346 ^~ reg307) ? ((8'haa) ? reg343 : wire324) : (!reg303)) ?
              $unsigned((~reg331)) : (reg317 ^~ reg300[(5'h12):(4'hd)])) : reg300[(4'h8):(3'h6)])))
        begin
          if (wire324[(3'h4):(1'h1)])
            begin
              reg401 = reg396;
              reg402 <= ($signed($signed($unsigned((-reg337)))) <= (reg365 ?
                  $signed($unsigned($unsigned((8'hb4)))) : $unsigned((!(reg372 ?
                      reg375 : reg339)))));
              reg403 <= $signed(reg346);
              reg404 <= wire293[(2'h2):(2'h2)];
            end
          else
            begin
              reg402 <= (~&(reg400 ?
                  reg300[(1'h1):(1'h0)] : (~^$unsigned((reg387 < reg387)))));
              reg403 <= (8'ha8);
            end
        end
      else
        begin
          if ({reg392})
            begin
              reg401 = (reg350[(2'h2):(2'h2)] & (8'hbb));
              reg405 = wire294[(1'h0):(1'h0)];
              reg406 = (~|(reg350 ? wire291 : reg397[(1'h0):(1'h0)]));
              reg407 <= reg335;
              reg408 <= {$signed($unsigned({(reg346 >> reg321), reg317})),
                  $unsigned($signed(((~&reg331) < wire295[(1'h0):(1'h0)])))};
            end
          else
            begin
              reg402 <= wire361[(2'h2):(1'h0)];
              reg405 = {(($unsigned({wire297,
                      reg303}) && $unsigned(reg365[(2'h2):(1'h1)])) >= ({(reg344 ?
                              reg363 : reg337),
                          (!reg300)} ?
                      ($unsigned(reg332) ?
                          $unsigned(reg408) : ((8'ha5) >= wire360)) : ((&forvar389) || (reg337 != reg353)))),
                  (^~{((reg317 != reg344) ?
                          $unsigned(reg331) : $signed(reg365)),
                      ({reg346, (7'h41)} ? $unsigned(reg400) : (+wire289))})};
              reg406 = reg354;
            end
          for (forvar409 = (1'h0); (forvar409 < (2'h3)); forvar409 = (forvar409 + (1'h1)))
            begin
              reg410 = (((((reg403 ^ wire360) & ((8'hb6) ?
                          (7'h44) : (8'had))) >>> $signed((reg408 <<< reg332))) ?
                      reg396[(2'h2):(1'h0)] : {$unsigned($unsigned(wire294)),
                          {reg317, $signed(forvar395)}}) ?
                  $signed({($unsigned(reg406) <= $unsigned(wire361)),
                      {(~^(8'had)),
                          (wire295 ?
                              wire293 : reg320)}}) : ((forvar409[(1'h1):(1'h0)] ?
                      $unsigned((reg332 << reg347)) : reg350) <= $signed(reg353[(2'h2):(2'h2)])));
              reg411 = reg402;
              reg412 = reg331;
            end
          reg413 = {$unsigned(reg337)};
          if (wire296)
            begin
              reg414 <= (wire291 + (~(reg403[(3'h6):(3'h5)] - ((wire294 >> reg302) != (reg353 >> wire294)))));
              reg415 <= reg303;
              reg416 = wire290;
              reg417 = (($unsigned($signed((8'hbe))) ?
                  (~^$unsigned((^reg307))) : reg343) != reg318[(1'h1):(1'h0)]);
              reg418 <= ((^$unsigned($unsigned($unsigned(wire293)))) < reg401);
            end
          else
            begin
              reg416 = {(-forvar388),
                  ((^~($signed(reg300) ?
                      $signed(reg317) : $unsigned(reg417))) >= reg323)};
              reg418 <= $signed({reg343});
              reg419 = (reg335 ?
                  $signed($signed(((reg307 ? reg368 : reg375) ?
                      reg344 : {reg397}))) : $unsigned((reg372 < ((reg407 | reg309) >= reg318))));
            end
        end
    end
  assign wire420 = (({reg377} == (7'h40)) ?
                       (!($signed((reg314 ? wire289 : reg320)) ?
                           (~&(wire324 ?
                               reg337 : reg363)) : reg418[(4'hd):(4'hb)])) : reg335);
  always
    @(posedge clk) begin
      reg421 = (~^({reg391, wire293} ?
          (reg318 ?
              $unsigned($signed(reg331)) : reg390) : (+$signed((wire296 & wire295)))));
      reg422 = (($signed((((8'ha5) + reg350) > $signed(wire324))) ?
              (8'hae) : $signed((reg393 ?
                  $signed(reg321) : (reg332 & wire289)))) ?
          (+wire291) : $unsigned($unsigned({$signed(reg414),
              $signed(wire294)})));
      reg423 = reg343;
    end
  assign wire424 = wire293[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg425 = ((|$unsigned((~|$unsigned(wire295)))) | wire361);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module125
#(parameter param242 = ((^~((!(-(8'hb6))) <<< (((7'h41) >= (7'h42)) ? ((8'hae) ? (8'hae) : (8'h9e)) : (~|(8'hb7))))) ? (((((8'hb8) ? (8'ha3) : (8'ha5)) || {(8'hac)}) <= ((~|(7'h42)) ? ((8'haf) ? (7'h42) : (7'h40)) : (~|(7'h43)))) ? ((((8'hbd) < (8'hab)) ? (+(8'ha6)) : (^~(7'h41))) >= (((8'haa) ? (7'h41) : (8'hb0)) ? (+(8'haa)) : (~|(8'ha0)))) : (8'hb4)) : ({{((8'hba) ? (7'h42) : (8'ha7))}} * ({{(8'ha2), (8'ha4)}} ? ((8'hb7) ~^ ((8'hb4) ? (7'h43) : (8'hb7))) : (((8'hbd) ? (8'hb4) : (8'hbf)) <= ((8'haf) != (8'hac)))))))
(y, clk, wire129, wire128, wire127, wire126);
  output wire [(32'h625):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire129;
  input wire [(4'h8):(1'h0)] wire128;
  input wire signed [(4'h9):(1'h0)] wire127;
  input wire signed [(4'hb):(1'h0)] wire126;
  wire [(4'hc):(1'h0)] wire207;
  wire [(2'h3):(1'h0)] wire131;
  wire [(5'h12):(1'h0)] wire130;
  reg signed [(4'hc):(1'h0)] reg237 = (1'h0);
  reg [(2'h2):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg230 = (1'h0);
  reg [(4'hb):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg228 = (1'h0);
  reg [(4'ha):(1'h0)] reg227 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg217 = (1'h0);
  reg [(5'h18):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg211 = (1'h0);
  reg signed [(4'he):(1'h0)] reg208 = (1'h0);
  reg [(4'hb):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] reg202 = (1'h0);
  reg [(5'h12):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg190 = (1'h0);
  reg signed [(4'he):(1'h0)] reg188 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg185 = (1'h0);
  reg [(3'h6):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg175 = (1'h0);
  reg [(5'h17):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg163 = (1'h0);
  reg [(4'ha):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg159 = (1'h0);
  reg [(3'h5):(1'h0)] reg153 = (1'h0);
  reg [(3'h4):(1'h0)] reg151 = (1'h0);
  reg [(4'hd):(1'h0)] reg148 = (1'h0);
  reg [(4'hd):(1'h0)] reg147 = (1'h0);
  reg [(5'h14):(1'h0)] reg146 = (1'h0);
  reg [(4'hc):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg143 = (1'h0);
  reg [(4'h9):(1'h0)] reg138 = (1'h0);
  reg [(5'h12):(1'h0)] reg137 = (1'h0);
  reg [(3'h5):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg135 = (1'h0);
  reg [(5'h16):(1'h0)] reg133 = (1'h0);
  reg [(4'h9):(1'h0)] reg241 = (1'h0);
  reg [(5'h15):(1'h0)] reg240 = (1'h0);
  reg [(4'hc):(1'h0)] reg239 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg234 = (1'h0);
  reg [(4'h8):(1'h0)] reg233 = (1'h0);
  reg [(5'h16):(1'h0)] reg232 = (1'h0);
  reg [(4'ha):(1'h0)] reg226 = (1'h0);
  reg [(5'h16):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar224 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar219 = (1'h0);
  reg [(2'h2):(1'h0)] reg218 = (1'h0);
  reg [(4'ha):(1'h0)] reg223 = (1'h0);
  reg [(5'h18):(1'h0)] forvar222 = (1'h0);
  reg [(2'h3):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg219 = (1'h0);
  reg [(4'hb):(1'h0)] forvar218 = (1'h0);
  reg [(4'hc):(1'h0)] reg215 = (1'h0);
  reg signed [(4'he):(1'h0)] reg213 = (1'h0);
  reg [(5'h17):(1'h0)] reg212 = (1'h0);
  reg [(5'h17):(1'h0)] forvar208 = (1'h0);
  reg signed [(4'he):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg209 = (1'h0);
  reg signed [(4'he):(1'h0)] reg206 = (1'h0);
  reg [(5'h18):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg203 = (1'h0);
  reg [(5'h16):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg199 = (1'h0);
  reg [(4'ha):(1'h0)] forvar198 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar197 = (1'h0);
  reg [(4'h8):(1'h0)] reg196 = (1'h0);
  reg [(4'h8):(1'h0)] reg194 = (1'h0);
  reg [(3'h4):(1'h0)] forvar191 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg189 = (1'h0);
  reg [(5'h17):(1'h0)] reg187 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg186 = (1'h0);
  reg [(2'h2):(1'h0)] forvar184 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar183 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg181 = (1'h0);
  reg [(5'h16):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg177 = (1'h0);
  reg [(5'h14):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar170 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar168 = (1'h0);
  reg [(5'h12):(1'h0)] reg169 = (1'h0);
  reg [(3'h6):(1'h0)] reg168 = (1'h0);
  reg [(4'h9):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg166 = (1'h0);
  reg [(4'ha):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar162 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg158 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar156 = (1'h0);
  reg [(5'h11):(1'h0)] reg155 = (1'h0);
  reg [(3'h7):(1'h0)] reg154 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg152 = (1'h0);
  reg [(5'h18):(1'h0)] reg150 = (1'h0);
  reg [(3'h6):(1'h0)] reg149 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar132 = (1'h0);
  reg [(5'h14):(1'h0)] reg142 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg141 = (1'h0);
  reg [(5'h10):(1'h0)] forvar140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg139 = (1'h0);
  reg [(4'h8):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg132 = (1'h0);
  assign y = {wire207,
                 wire131,
                 wire130,
                 reg237,
                 reg235,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg217,
                 reg216,
                 reg214,
                 reg211,
                 reg208,
                 reg204,
                 reg202,
                 reg200,
                 reg195,
                 reg193,
                 reg192,
                 reg190,
                 reg188,
                 reg185,
                 reg178,
                 reg176,
                 reg175,
                 reg174,
                 reg172,
                 reg165,
                 reg163,
                 reg161,
                 reg159,
                 reg153,
                 reg151,
                 reg148,
                 reg147,
                 reg146,
                 reg144,
                 reg140,
                 reg143,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg133,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg236,
                 reg234,
                 reg233,
                 reg232,
                 reg226,
                 reg225,
                 forvar224,
                 forvar219,
                 reg218,
                 reg223,
                 forvar222,
                 reg221,
                 reg220,
                 reg219,
                 forvar218,
                 reg215,
                 reg213,
                 reg212,
                 forvar208,
                 reg210,
                 reg209,
                 reg206,
                 reg205,
                 reg203,
                 reg201,
                 reg199,
                 forvar198,
                 forvar197,
                 reg196,
                 reg194,
                 forvar191,
                 reg189,
                 reg187,
                 reg186,
                 forvar184,
                 forvar183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg177,
                 reg173,
                 reg171,
                 forvar170,
                 forvar168,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg164,
                 forvar162,
                 reg160,
                 reg158,
                 reg157,
                 forvar156,
                 reg155,
                 reg154,
                 reg152,
                 reg150,
                 reg149,
                 reg145,
                 forvar132,
                 reg142,
                 reg141,
                 forvar140,
                 reg139,
                 reg134,
                 reg132,
                 (1'h0)};
  assign wire130 = wire126;
  assign wire131 = (wire129[(1'h0):(1'h0)] && (wire126[(4'h9):(2'h3)] ?
                       ({wire127[(2'h2):(1'h0)]} << (wire129 >>> (&(8'hba)))) : wire126[(4'h9):(3'h4)]));
  always
    @(posedge clk) begin
      if (((({wire131, wire131} ?
              ($signed(wire127) < (wire128 ?
                  wire129 : (7'h47))) : wire127[(3'h7):(1'h1)]) ?
          ($signed((wire128 ? wire127 : wire129)) || ($signed(wire127) ?
              (wire128 >= (8'hb9)) : $signed(wire129))) : (wire127[(3'h7):(3'h5)] ?
              {(wire126 | wire130)} : $signed($signed(wire130)))) ~^ wire130[(4'hc):(1'h1)]))
        begin
          reg132 = $signed(((({wire126} ?
              (wire129 ? wire128 : wire129) : {wire128,
                  wire130}) | (^~wire130[(2'h2):(1'h0)])) < (&wire128[(2'h2):(2'h2)])));
          reg133 <= ((wire126[(2'h2):(1'h1)] || $signed({(+wire128)})) ?
              (wire127 <<< wire131[(1'h0):(1'h0)]) : {(&(~^(reg132 ?
                      wire128 : wire126))),
                  (8'hb7)});
          if ($unsigned(wire126[(4'h8):(1'h0)]))
            begin
              reg134 = ((-(~^((~&wire131) > (wire131 ? wire128 : wire127)))) ?
                  wire129[(2'h2):(1'h1)] : {reg132});
            end
          else
            begin
              reg135 <= ($signed({{(!wire127)}}) <<< ((wire129[(2'h3):(1'h0)] != $unsigned({reg134})) ?
                  wire130 : wire127));
              reg136 <= ({($signed($unsigned(reg132)) && $signed((reg134 == wire129)))} ?
                  $signed(reg133[(4'hc):(2'h3)]) : wire131[(2'h3):(2'h2)]);
              reg137 <= (((($signed(reg136) <= (8'ha1)) || $signed($signed(reg136))) - $unsigned(reg136)) <<< (reg135 ?
                  $signed($signed((8'h9d))) : (reg135 ? wire126 : reg134)));
              reg138 <= $signed(({wire128,
                  (^~(reg134 ?
                      reg137 : wire131))} - $signed((reg136[(2'h3):(1'h1)] ?
                  {wire126} : (~^wire129)))));
              reg139 = reg137;
            end
          for (forvar140 = (1'h0); (forvar140 < (1'h1)); forvar140 = (forvar140 + (1'h1)))
            begin
              reg141 = (~|(^~($signed({reg132, reg135}) ?
                  wire130 : $signed((~reg138)))));
              reg142 = ((8'ha0) ?
                  $unsigned($signed({((8'hb3) || reg141)})) : (~|(^~wire130)));
              reg143 <= reg139[(2'h3):(2'h3)];
            end
        end
      else
        begin
          for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg134 = ($unsigned(((reg141 ? (!wire128) : (|(8'hb5))) ?
                  reg143[(4'ha):(3'h6)] : reg134[(2'h3):(1'h0)])) >= wire130);
              reg135 <= $signed({$unsigned(($unsigned(forvar140) ?
                      (~(8'hb8)) : $unsigned(wire130)))});
            end
          reg139 = wire127[(4'h8):(3'h7)];
          if ((~^((|$unsigned((reg143 == reg133))) ?
              reg141[(3'h6):(1'h0)] : (((forvar132 & reg133) ?
                      (reg142 ? reg132 : wire128) : (7'h49)) ?
                  $signed($signed(reg141)) : $signed(wire131)))))
            begin
              reg140 <= (~|(~(({reg139, reg143} ?
                  reg134 : (^~wire128)) - (^~wire131))));
              reg143 <= {wire127, wire131[(2'h3):(2'h3)]};
            end
          else
            begin
              reg141 = $unsigned($unsigned({$signed(reg133)}));
            end
          reg144 <= $unsigned($signed(reg140[(4'he):(4'hc)]));
          reg145 = reg143;
        end
      reg146 <= $signed((8'hb1));
      reg147 <= {reg136[(1'h0):(1'h0)],
          $unsigned($signed((wire128 || $unsigned(wire130))))};
      reg148 <= (reg141[(2'h3):(2'h3)] ?
          $signed((~^({wire127, reg135} && (reg147 ?
              reg133 : reg141)))) : wire127);
      reg149 = reg147;
    end
  always
    @(posedge clk) begin
      if ((((+$unsigned($unsigned(wire127))) ?
              (($signed(reg140) << reg148) ~^ reg137) : ((+{reg146}) ?
                  ($unsigned(wire129) - $unsigned((8'ha5))) : reg143)) ?
          (&$signed($unsigned($signed(reg146)))) : wire129))
        begin
          if ($unsigned(($signed(((reg133 ? wire128 : reg135) ?
              (reg148 <<< wire127) : $unsigned(reg144))) >>> reg136[(2'h3):(1'h0)])))
            begin
              reg150 = $signed(reg140[(5'h14):(4'h9)]);
              reg151 <= (7'h41);
            end
          else
            begin
              reg151 <= ($signed(reg138) ?
                  (+$signed((wire130[(5'h11):(4'hb)] - $signed(reg143)))) : ((reg151 ?
                          ((|wire130) ?
                              (reg137 >= (8'hbc)) : reg138) : $signed((reg144 ?
                              (8'hb5) : reg133))) ?
                      (-({reg147} == (reg136 <<< reg151))) : {(^$unsigned(wire128))}));
              reg152 = (~&$signed(((~$signed(wire131)) ?
                  reg148 : ({wire129} > wire127[(2'h2):(1'h0)]))));
              reg153 <= {(((~(reg144 - (7'h42))) || reg136[(2'h3):(2'h3)]) >> $signed(reg143))};
              reg154 = wire130[(1'h0):(1'h0)];
              reg155 = ((+(|$unsigned((reg137 | reg135)))) ?
                  (reg150[(5'h11):(3'h6)] ^~ reg147) : ($signed($signed(wire127[(3'h4):(2'h2)])) ~^ reg138[(3'h6):(2'h2)]));
            end
          for (forvar156 = (1'h0); (forvar156 < (1'h0)); forvar156 = (forvar156 + (1'h1)))
            begin
              reg157 = (wire129 || (8'h9f));
              reg158 = wire126[(3'h5):(2'h2)];
            end
          reg159 <= $signed((!(^$signed(wire129[(3'h4):(2'h3)]))));
          reg160 = ($unsigned(reg133[(5'h10):(3'h5)]) ^ $signed({((reg144 ?
                      reg135 : (8'h9e)) ?
                  (8'hb5) : $unsigned((7'h45))),
              $signed(reg148)}));
        end
      else
        begin
          reg151 <= {reg155[(4'h8):(2'h2)],
              (~|$unsigned(forvar156[(3'h6):(3'h4)]))};
        end
      reg161 <= (&wire126);
      for (forvar162 = (1'h0); (forvar162 < (1'h0)); forvar162 = (forvar162 + (1'h1)))
        begin
          reg163 <= reg135[(2'h2):(1'h0)];
          reg164 = reg147[(3'h5):(2'h3)];
          reg165 <= (7'h41);
        end
    end
  always
    @(posedge clk) begin
      reg166 = $unsigned(reg138[(4'h9):(2'h3)]);
      reg167 = reg135;
    end
  always
    @(posedge clk) begin
      if (($unsigned((~reg133[(5'h13):(3'h7)])) >> $signed($signed((reg144 != (reg159 << reg146))))))
        begin
          reg168 = wire131[(1'h1):(1'h0)];
          reg169 = reg138[(1'h1):(1'h1)];
        end
      else
        begin
          for (forvar168 = (1'h0); (forvar168 < (2'h2)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 = $signed((~reg137[(4'hb):(3'h6)]));
            end
          for (forvar170 = (1'h0); (forvar170 < (2'h2)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 = ({reg165[(5'h11):(3'h4)]} << forvar168[(4'h9):(2'h3)]);
              reg172 <= {wire126[(3'h5):(2'h3)], reg144};
              reg173 = (((($unsigned(reg153) - reg135[(3'h4):(1'h1)]) < $unsigned((7'h44))) ~^ reg146[(3'h6):(1'h1)]) ?
                  $signed((-((reg161 ~^ wire127) ?
                      $signed(reg138) : reg135[(3'h6):(2'h2)]))) : (-$signed($unsigned($signed(wire127)))));
              reg174 <= $signed(wire131[(1'h1):(1'h1)]);
              reg175 <= $unsigned(reg148[(4'ha):(4'ha)]);
            end
          if (($unsigned(reg174[(5'h17):(5'h12)]) ?
              reg173[(3'h4):(2'h3)] : (~^reg171)))
            begin
              reg176 <= reg148[(2'h3):(2'h3)];
              reg177 = forvar170[(2'h2):(1'h1)];
              reg178 <= {(^~wire126)};
              reg179 = $signed($signed(((reg146 ?
                  (reg159 << reg143) : reg144[(4'h8):(1'h0)]) ^ $signed(reg151[(2'h3):(2'h3)]))));
              reg180 = $signed(reg144);
            end
          else
            begin
              reg176 <= $signed((!(^$signed((reg161 ? forvar168 : reg140)))));
            end
          reg181 = ((~reg153) ?
              (reg137[(4'hb):(2'h3)] ?
                  ((^(&reg140)) ?
                      ((|reg144) ?
                          (reg180 >= reg137) : reg173) : $signed((~^reg148))) : ((reg151 ?
                      wire127 : {reg168,
                          reg147}) << ($signed((7'h47)) || {(8'hb2)}))) : reg151[(2'h2):(2'h2)]);
        end
      reg182 = (^~((!reg163) + $signed(reg136[(3'h4):(2'h2)])));
      for (forvar183 = (1'h0); (forvar183 < (3'h4)); forvar183 = (forvar183 + (1'h1)))
        begin
          for (forvar184 = (1'h0); (forvar184 < (3'h4)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 <= ((-$unsigned($signed({(8'hab)}))) ^ (($unsigned($signed((7'h41))) << $signed(reg169[(4'h8):(3'h6)])) ?
                  reg177 : $signed(((!reg133) || {reg138, reg144}))));
              reg186 = (~&reg135[(4'hb):(4'ha)]);
              reg187 = reg182[(1'h0):(1'h0)];
              reg188 <= {reg178[(1'h1):(1'h1)]};
            end
          if ($signed((~&forvar184)))
            begin
              reg189 = $unsigned(($signed(($unsigned(wire126) <<< $unsigned((8'ha0)))) < (8'ha5)));
            end
          else
            begin
              reg189 = forvar184[(1'h1):(1'h0)];
              reg190 <= ((reg133 ?
                      reg187[(3'h7):(2'h2)] : (($unsigned(reg151) <<< $unsigned(reg169)) ?
                          (reg180 >>> {reg175, (8'hbc)}) : (~(reg171 ?
                              reg171 : reg179)))) ?
                  $unsigned(($signed((8'hb3)) ?
                      {(8'ha9),
                          $unsigned((8'hb3))} : (|$unsigned(wire129)))) : $signed($unsigned(((reg181 & forvar183) ?
                      wire129[(1'h1):(1'h0)] : reg151[(3'h4):(1'h0)]))));
            end
          for (forvar191 = (1'h0); (forvar191 < (1'h0)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= reg138;
              reg193 <= $unsigned(reg133);
              reg194 = ((8'hb4) ?
                  $unsigned({$signed((reg133 >> reg172)),
                      reg174[(5'h16):(5'h14)]}) : reg181);
              reg195 <= (~$signed($signed($signed((reg148 || (8'ha4))))));
              reg196 = ($signed({($unsigned((7'h40)) <= (wire130 ?
                      reg165 : (8'ha6)))}) != ({(reg194 ?
                          wire127 : (reg136 ? (7'h47) : reg177)),
                      ((forvar191 + (8'hbd)) ?
                          (!(8'ha0)) : $unsigned(reg174))} ?
                  reg168 : ((~reg143[(5'h13):(4'h8)]) ?
                      $signed(reg178[(1'h0):(1'h0)]) : (~|$signed(reg178)))));
            end
        end
      for (forvar197 = (1'h0); (forvar197 < (1'h1)); forvar197 = (forvar197 + (1'h1)))
        begin
          for (forvar198 = (1'h0); (forvar198 < (1'h0)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 = $unsigned((~&(|{$signed(reg180)})));
              reg200 <= (reg179 ?
                  ($signed($unsigned($signed(wire128))) != $signed($unsigned(wire127))) : reg161[(1'h0):(1'h0)]);
              reg201 = (~$signed(reg194[(1'h1):(1'h0)]));
              reg202 <= (reg195 & {reg196});
              reg203 = $signed({{{$signed(reg163),
                          (reg179 ? wire128 : reg174)}}});
            end
          if ((($signed((!(8'haa))) <<< ($unsigned($unsigned(reg187)) | (|forvar191[(1'h1):(1'h0)]))) == reg200))
            begin
              reg204 <= reg165[(3'h6):(2'h3)];
              reg205 = ((($signed(reg187) <= (|(reg133 < reg133))) && reg135) || $unsigned((~&$signed($unsigned(reg202)))));
              reg206 = forvar170[(1'h1):(1'h1)];
            end
          else
            begin
              reg204 <= reg194;
              reg205 = reg187[(4'hf):(2'h2)];
              reg206 = {({(reg205[(1'h1):(1'h0)] == $unsigned(reg202))} != wire128[(1'h1):(1'h1)]),
                  (reg171[(3'h5):(1'h1)] ?
                      (+{$signed((8'ha9)),
                          reg176[(4'hb):(4'hb)]}) : ($unsigned($signed(reg169)) | reg186))};
            end
        end
    end
  assign wire207 = $unsigned(((!$signed(reg165[(3'h7):(3'h4)])) ?
                       $unsigned(((reg133 ?
                           reg136 : reg146) ^ $unsigned(reg192))) : (reg151[(1'h0):(1'h0)] ?
                           $signed($unsigned(reg143)) : $signed($unsigned(reg137)))));
  always
    @(posedge clk) begin
      if ($unsigned((-((^~(reg140 ?
          reg200 : reg192)) <= reg195[(3'h5):(1'h1)]))))
        begin
          if (reg188)
            begin
              reg208 <= $signed({{(reg147 + reg151[(1'h1):(1'h1)]),
                      $unsigned(reg144)},
                  (((reg175 ? reg133 : reg192) ?
                          reg137[(4'ha):(4'h9)] : (reg137 << reg138)) ?
                      (8'hb4) : ((reg136 ? reg137 : wire127) ^ (reg163 ?
                          wire127 : reg161)))});
            end
          else
            begin
              reg209 = {(reg185 ?
                      (((reg135 ? reg193 : (8'ha5)) ?
                          (~^wire131) : reg159[(4'h8):(2'h2)]) <<< (^~$unsigned(reg138))) : (~$unsigned((+reg136)))),
                  wire129};
              reg210 = (|((reg146[(2'h3):(2'h2)] ?
                      (|$signed(reg133)) : ((^~reg209) ?
                          (reg202 ^~ reg136) : reg176)) ?
                  wire131 : $unsigned(reg151)));
            end
        end
      else
        begin
          for (forvar208 = (1'h0); (forvar208 < (2'h2)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg211 <= (+reg153);
              reg212 = $signed({(~|(!$unsigned(wire129))), $signed(reg148)});
            end
          reg213 = $unsigned(reg144[(1'h1):(1'h0)]);
          reg214 <= (reg133 ?
              ((~&({reg190, wire127} ?
                  (!reg138) : reg213)) && ((reg195[(2'h2):(1'h0)] << wire130) ?
                  (~^reg176) : $unsigned(reg159))) : $signed(reg178));
        end
    end
  always
    @(posedge clk) begin
      if (((~&(wire207 ? $signed($signed(reg204)) : {(reg153 ~^ wire130)})) ?
          reg136[(1'h1):(1'h0)] : {(~|{$signed(reg211)}),
              $unsigned(($unsigned(reg174) ?
                  $unsigned(reg163) : (wire131 ? wire129 : reg165)))}))
        begin
          reg215 = ((reg137[(1'h0):(1'h0)] ?
                  ({((8'ha9) ? reg165 : (7'h46)), (8'hbd)} ?
                      {(reg188 ? reg204 : reg137),
                          $signed(wire207)} : $signed((reg163 ?
                          reg195 : reg165))) : (reg174 + ($unsigned(reg174) & (-reg147)))) ?
              (&(wire127[(3'h6):(1'h1)] ?
                  {reg185, (^~reg135)} : ({reg190} * (reg200 ?
                      (8'ha2) : (7'h40))))) : $unsigned(reg172[(4'h9):(3'h4)]));
          reg216 <= (8'ha8);
          reg217 <= wire129;
          for (forvar218 = (1'h0); (forvar218 < (2'h2)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 = $unsigned((($signed((reg165 ? wire130 : (8'hb3))) ?
                  $unsigned(wire131) : $unsigned((~|(8'hb5)))) > ($unsigned(reg172) ?
                  reg202 : $signed({reg138}))));
              reg220 = (|reg148[(2'h3):(2'h3)]);
              reg221 = (reg143 ?
                  $unsigned({$signed(reg195),
                      reg185[(2'h2):(1'h0)]}) : (7'h42));
            end
          for (forvar222 = (1'h0); (forvar222 < (2'h3)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 = (^reg159[(4'hc):(4'hc)]);
            end
        end
      else
        begin
          reg216 <= {reg136[(1'h0):(1'h0)],
              ((({reg185} > (reg133 || reg193)) != reg216) & $unsigned(reg163))};
          reg218 = (forvar218[(2'h2):(1'h1)] | $unsigned(reg146));
          for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 = (!$unsigned(((+{reg163, reg220}) ?
                  (+(reg165 != wire129)) : $signed(((7'h4a) ^ reg192)))));
            end
        end
      for (forvar224 = (1'h0); (forvar224 < (2'h3)); forvar224 = (forvar224 + (1'h1)))
        begin
          if ((reg140[(4'hb):(3'h6)] >> {$unsigned($unsigned(reg217))}))
            begin
              reg225 = reg178[(1'h1):(1'h0)];
              reg226 = (&reg175);
              reg227 <= $signed(wire130[(4'hc):(2'h3)]);
            end
          else
            begin
              reg227 <= (7'h43);
              reg228 <= (wire129[(3'h4):(2'h3)] > ((|reg204) ^ $signed($unsigned(wire128))));
              reg229 <= $signed(((~^$unsigned(reg193[(4'ha):(3'h7)])) ?
                  (8'hb2) : reg193[(4'h8):(3'h4)]));
              reg230 <= (+($unsigned((+reg192[(4'he):(4'hc)])) ?
                  {($signed((8'hbb)) ^ (reg174 ?
                          reg216 : reg214))} : $unsigned(forvar224[(3'h5):(1'h1)])));
              reg231 <= $unsigned(((~&((reg218 | wire130) ?
                      (reg217 || reg172) : $signed(reg218))) ?
                  {reg140,
                      $unsigned((reg221 ?
                          reg193 : reg135))} : ($signed((reg215 - reg148)) ?
                      {reg220} : ((reg192 < reg193) ?
                          reg136[(1'h1):(1'h0)] : reg144[(1'h1):(1'h1)]))));
            end
          if ({$signed($signed((reg136 ? {reg230} : wire131))),
              ((wire207 ? reg218[(1'h0):(1'h0)] : $signed($unsigned(reg148))) ?
                  reg218[(1'h1):(1'h1)] : $unsigned($signed(wire131[(1'h0):(1'h0)])))})
            begin
              reg232 = reg159[(5'h10):(1'h1)];
              reg233 = reg172[(5'h13):(4'hb)];
              reg234 = ($signed((|(reg175[(5'h11):(5'h11)] != (wire130 & reg192)))) >> wire207[(4'hc):(4'hb)]);
              reg235 <= {((($unsigned(wire126) != (~^reg227)) ?
                          (~|reg135) : $signed(((7'h4a) ? reg151 : reg143))) ?
                      wire127[(3'h7):(2'h2)] : $signed(({reg175} & $unsigned(forvar219))))};
            end
          else
            begin
              reg232 = reg136[(1'h1):(1'h0)];
              reg233 = (((7'h48) ? reg147 : $unsigned($signed(wire207))) ?
                  $unsigned((({(8'haa)} & reg148) + (wire131[(1'h0):(1'h0)] >>> reg192[(4'hb):(4'h9)]))) : $signed(reg217));
              reg234 = reg172;
            end
          if (forvar218)
            begin
              reg236 = $signed((reg233 ?
                  ((8'ha5) ?
                      $unsigned((~|wire127)) : (reg228 >> $unsigned(wire207))) : (~^$signed((reg147 ?
                      reg231 : reg163)))));
              reg237 <= wire130[(5'h11):(5'h10)];
            end
          else
            begin
              reg237 <= (~&reg161[(3'h5):(2'h2)]);
              reg238 = (~^$signed($unsigned((~$signed((8'ha0))))));
              reg239 = reg172[(3'h6):(1'h1)];
              reg240 = reg232[(3'h4):(1'h0)];
              reg241 = reg148[(3'h5):(3'h5)];
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module803  (y, clk, wire807, wire806, wire805, wire804);
  output wire [(32'hfe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire807;
  input wire signed [(5'h10):(1'h0)] wire806;
  input wire [(3'h7):(1'h0)] wire805;
  input wire signed [(3'h7):(1'h0)] wire804;
  wire signed [(5'h12):(1'h0)] wire822;
  wire signed [(4'ha):(1'h0)] wire821;
  wire signed [(5'h17):(1'h0)] wire820;
  wire signed [(4'hd):(1'h0)] wire819;
  wire [(5'h11):(1'h0)] wire817;
  wire [(5'h18):(1'h0)] wire816;
  wire signed [(4'he):(1'h0)] wire815;
  wire signed [(3'h6):(1'h0)] wire811;
  wire [(5'h15):(1'h0)] wire810;
  wire signed [(5'h11):(1'h0)] wire809;
  wire signed [(2'h2):(1'h0)] wire808;
  reg [(5'h18):(1'h0)] reg823 = (1'h0);
  reg [(3'h7):(1'h0)] reg812 = (1'h0);
  reg [(5'h15):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg818 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg814 = (1'h0);
  reg [(4'hc):(1'h0)] reg813 = (1'h0);
  assign y = {wire822,
                 wire821,
                 wire820,
                 wire819,
                 wire817,
                 wire816,
                 wire815,
                 wire811,
                 wire810,
                 wire809,
                 wire808,
                 reg823,
                 reg812,
                 reg824,
                 reg818,
                 reg814,
                 reg813,
                 (1'h0)};
  assign wire808 = (wire807[(3'h7):(3'h7)] ?
                       wire804[(3'h4):(2'h2)] : wire806[(3'h5):(3'h5)]);
  assign wire809 = wire804[(3'h4):(2'h2)];
  assign wire810 = wire809;
  assign wire811 = (+(8'ha2));
  always
    @(posedge clk) begin
      reg812 <= ((8'h9d) ?
          (8'ha3) : ((~^($signed(wire811) ?
                  wire807[(4'hc):(2'h3)] : $signed((8'haa)))) ?
              wire810[(5'h10):(4'h8)] : (($signed(wire810) | wire811) ?
                  $signed(wire811) : $signed({wire809, wire806}))));
      reg813 = reg812;
      reg814 = $unsigned(((wire807[(3'h4):(3'h4)] ?
          wire807 : ((^~reg813) ?
              $unsigned((8'ha7)) : $unsigned(reg812))) + (-((+wire807) ~^ (|wire808)))));
    end
  assign wire815 = (&wire807[(3'h5):(1'h0)]);
  assign wire816 = $signed(($unsigned(((8'hac) ?
                       wire809[(2'h3):(1'h0)] : (wire810 != wire806))) >> (wire810 < ($unsigned(wire808) != reg812))));
  assign wire817 = wire808[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg818 = $unsigned($signed(({wire806, wire804} >= ({wire805,
          wire815} ^~ (8'hb9)))));
    end
  assign wire819 = wire815;
  assign wire820 = wire808;
  assign wire821 = ({wire804[(1'h0):(1'h0)]} ?
                       wire806[(2'h3):(1'h1)] : (8'hb2));
  assign wire822 = (~$signed(((wire811 ?
                           ((8'ha7) < wire810) : $unsigned(reg812)) ?
                       (!(reg812 ? wire821 : wire816)) : {$signed(wire816),
                           wire820})));
  always
    @(posedge clk) begin
      reg823 <= wire821;
      reg824 = (($unsigned($unsigned($unsigned(wire819))) && ($signed((wire820 ?
              wire819 : wire811)) | (8'haa))) ?
          wire806[(2'h2):(2'h2)] : $unsigned(wire820));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module705
#(parameter param799 = {(!((((8'ha0) < (8'hab)) != (-(7'h40))) ~^ (^~((8'h9e) < (8'had))))), (((((8'h9f) | (8'hb1)) || ((7'h45) >> (8'ha2))) ? {((8'hae) >> (8'h9f))} : (((8'ha6) ? (8'ha9) : (8'ha7)) ? (~^(7'h42)) : ((8'hb4) ? (8'hb1) : (8'had)))) ? (({(8'hbd), (8'ha9)} ? ((8'h9d) - (7'h49)) : {(8'hae)}) ? ({(8'hb8), (7'h48)} | (+(8'hae))) : {(-(8'hb3))}) : {(((7'h47) ? (8'h9d) : (8'hba)) < ((7'h45) ? (8'hb6) : (8'hb0)))})})
(y, clk, wire709, wire708, wire707, wire706);
  output wire [(32'h4c1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire709;
  input wire signed [(5'h10):(1'h0)] wire708;
  input wire signed [(5'h18):(1'h0)] wire707;
  input wire [(3'h5):(1'h0)] wire706;
  wire [(4'hb):(1'h0)] wire798;
  wire [(4'hb):(1'h0)] wire797;
  wire signed [(4'he):(1'h0)] wire769;
  wire signed [(5'h12):(1'h0)] wire761;
  wire signed [(4'h9):(1'h0)] wire760;
  wire signed [(5'h13):(1'h0)] wire759;
  wire signed [(4'he):(1'h0)] wire733;
  wire [(5'h17):(1'h0)] wire732;
  wire signed [(5'h17):(1'h0)] wire731;
  wire signed [(5'h10):(1'h0)] wire730;
  wire signed [(4'hb):(1'h0)] wire729;
  wire [(5'h15):(1'h0)] wire714;
  wire signed [(4'hb):(1'h0)] wire713;
  wire [(3'h6):(1'h0)] wire712;
  wire signed [(3'h5):(1'h0)] wire711;
  wire [(3'h4):(1'h0)] wire710;
  reg [(4'hc):(1'h0)] reg796 = (1'h0);
  reg [(5'h18):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg792 = (1'h0);
  reg [(4'h8):(1'h0)] reg791 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg784 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg778 = (1'h0);
  reg [(3'h7):(1'h0)] reg777 = (1'h0);
  reg [(5'h16):(1'h0)] reg775 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg774 = (1'h0);
  reg [(4'hf):(1'h0)] reg773 = (1'h0);
  reg [(3'h6):(1'h0)] reg772 = (1'h0);
  reg [(4'ha):(1'h0)] reg771 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg767 = (1'h0);
  reg [(2'h2):(1'h0)] reg766 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg765 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg764 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg757 = (1'h0);
  reg [(4'hb):(1'h0)] reg756 = (1'h0);
  reg [(5'h18):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg750 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg747 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg745 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg742 = (1'h0);
  reg [(5'h12):(1'h0)] reg740 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg738 = (1'h0);
  reg [(4'he):(1'h0)] reg736 = (1'h0);
  reg [(5'h12):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg724 = (1'h0);
  reg [(5'h14):(1'h0)] reg722 = (1'h0);
  reg [(2'h2):(1'h0)] reg719 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg717 = (1'h0);
  reg [(4'hb):(1'h0)] reg716 = (1'h0);
  reg [(4'h8):(1'h0)] reg794 = (1'h0);
  reg [(5'h11):(1'h0)] forvar793 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg790 = (1'h0);
  reg [(2'h3):(1'h0)] reg789 = (1'h0);
  reg [(2'h2):(1'h0)] reg788 = (1'h0);
  reg [(4'hd):(1'h0)] reg787 = (1'h0);
  reg [(5'h16):(1'h0)] reg786 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg785 = (1'h0);
  reg [(5'h15):(1'h0)] forvar783 = (1'h0);
  reg [(4'hf):(1'h0)] reg782 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg781 = (1'h0);
  reg [(4'hb):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar779 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar776 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar771 = (1'h0);
  reg [(5'h10):(1'h0)] reg768 = (1'h0);
  reg [(4'hf):(1'h0)] forvar763 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg758 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg755 = (1'h0);
  reg [(5'h13):(1'h0)] reg753 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg752 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg751 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg748 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg746 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar744 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg739 = (1'h0);
  reg [(4'hb):(1'h0)] reg737 = (1'h0);
  reg [(5'h15):(1'h0)] forvar735 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar734 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar726 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg723 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar721 = (1'h0);
  reg [(2'h3):(1'h0)] reg720 = (1'h0);
  reg signed [(4'he):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg715 = (1'h0);
  assign y = {wire798,
                 wire797,
                 wire769,
                 wire761,
                 wire760,
                 wire759,
                 wire733,
                 wire732,
                 wire731,
                 wire730,
                 wire729,
                 wire714,
                 wire713,
                 wire712,
                 wire711,
                 wire710,
                 reg796,
                 reg795,
                 reg792,
                 reg791,
                 reg784,
                 reg778,
                 reg777,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg767,
                 reg766,
                 reg765,
                 reg764,
                 reg757,
                 reg756,
                 reg754,
                 reg750,
                 reg747,
                 reg745,
                 reg742,
                 reg740,
                 reg738,
                 reg736,
                 reg728,
                 reg725,
                 reg724,
                 reg722,
                 reg719,
                 reg717,
                 reg716,
                 reg794,
                 forvar793,
                 reg790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 forvar783,
                 reg782,
                 reg781,
                 reg780,
                 forvar779,
                 forvar776,
                 forvar771,
                 reg768,
                 forvar763,
                 reg762,
                 reg758,
                 reg755,
                 reg753,
                 reg752,
                 reg751,
                 forvar749,
                 reg748,
                 reg746,
                 forvar744,
                 forvar743,
                 reg741,
                 reg739,
                 reg737,
                 forvar735,
                 forvar734,
                 reg727,
                 forvar726,
                 reg723,
                 forvar721,
                 reg720,
                 reg718,
                 reg715,
                 (1'h0)};
  assign wire710 = wire706;
  assign wire711 = ($signed($unsigned(({wire706} <<< wire706[(2'h2):(1'h0)]))) != (^$unsigned(wire710[(1'h0):(1'h0)])));
  assign wire712 = (($signed($signed($unsigned(wire710))) ?
                           {wire709} : $signed((|{wire709}))) ?
                       $unsigned((~^wire706[(1'h1):(1'h1)])) : (($unsigned((wire707 ?
                           wire709 : wire708)) + ($unsigned(wire709) ?
                           (~&wire709) : wire708)) >= wire710));
  assign wire713 = ($unsigned((~|(^~wire706))) << {$signed(wire708), wire710});
  assign wire714 = ((wire708 & {((^~wire710) | $signed(wire707)),
                       wire707}) | $signed((((^(8'ha8)) ?
                           $signed(wire712) : {wire712, wire707}) ?
                       (wire713[(3'h6):(1'h0)] ?
                           wire706[(2'h3):(2'h3)] : {wire707}) : (^~(wire712 ?
                           wire709 : wire711)))));
  always
    @(posedge clk) begin
      if ((~^($unsigned({$unsigned(wire714)}) ?
          (((wire706 ?
              (7'h48) : wire714) ^ wire712) > (wire714 >> (wire707 && wire714))) : $signed((8'hb1)))))
        begin
          reg715 = ((8'hb3) + $unsigned(((^wire712[(2'h2):(1'h0)]) >>> $signed($signed((7'h40))))));
          reg716 <= wire711;
          reg717 <= ($signed((~&($unsigned(wire706) * (reg715 ?
                  reg715 : reg715)))) ?
              wire712[(3'h5):(2'h3)] : wire709[(5'h13):(5'h12)]);
          reg718 = wire713[(3'h4):(2'h3)];
          reg719 <= $unsigned($unsigned({((wire709 > reg718) ~^ $unsigned(reg716))}));
        end
      else
        begin
          reg715 = {$signed($signed(wire707))};
          if ((wire707 + (((~wire712) ?
                  reg716 : {wire712[(1'h0):(1'h0)],
                      (wire709 ? reg719 : (8'haa))}) ?
              {($unsigned(wire712) <<< wire714[(4'h8):(3'h4)])} : {{(^wire714)},
                  ($unsigned((8'hbe)) ? (~^wire712) : ((8'ha4) <= wire709))})))
            begin
              reg716 <= reg716;
              reg717 <= $unsigned(reg716);
              reg718 = (reg717[(3'h4):(1'h1)] ?
                  $unsigned($unsigned($signed($unsigned(wire714)))) : (~&($unsigned((!wire709)) ?
                      (&$unsigned(reg717)) : $signed((reg718 == wire712)))));
              reg719 <= ({(^~(wire706[(1'h0):(1'h0)] > $signed(reg715)))} >> ((reg717[(5'h13):(4'hf)] ?
                      ((wire711 ?
                          wire713 : wire709) < (~^(8'hb6))) : wire710[(1'h0):(1'h0)]) ?
                  reg715[(1'h1):(1'h0)] : wire712));
            end
          else
            begin
              reg718 = reg715[(1'h1):(1'h0)];
              reg719 <= ($signed((($unsigned(wire708) != (wire710 * reg718)) ?
                      $unsigned($unsigned(wire707)) : ($unsigned(reg716) ?
                          $signed(reg718) : {reg718}))) ?
                  (+($signed($unsigned(wire711)) ?
                      wire706 : ((-wire710) ?
                          (reg719 ^~ wire711) : wire708[(2'h2):(1'h1)]))) : (({wire707[(5'h15):(4'he)]} ?
                      $signed({wire708, reg719}) : {wire708[(3'h5):(2'h2)],
                          reg718[(4'hd):(4'hb)]}) == wire709));
              reg720 = (((&$unsigned(wire713)) ?
                      (~$signed(reg718[(4'h8):(3'h6)])) : (-((reg717 <<< reg718) <= wire714[(3'h5):(3'h4)]))) ?
                  ((^~($signed(reg717) ?
                          (wire713 ? reg719 : reg715) : (wire707 ?
                              (8'hb2) : wire714))) ?
                      (reg715[(1'h0):(1'h0)] ?
                          (reg717[(3'h6):(1'h1)] ^~ (wire710 <<< wire708)) : wire708) : $signed(((8'hb0) ?
                          ((8'hae) ^ wire706) : {wire713, reg716}))) : wire711);
            end
        end
      for (forvar721 = (1'h0); (forvar721 < (2'h2)); forvar721 = (forvar721 + (1'h1)))
        begin
          if ((7'h45))
            begin
              reg722 <= (!($signed(reg716[(4'h9):(2'h2)]) ?
                  reg719[(1'h1):(1'h0)] : $signed({$unsigned((8'hbf)),
                      (reg720 ? reg717 : wire707)})));
            end
          else
            begin
              reg723 = ($unsigned({reg717[(5'h15):(4'h9)],
                  ($signed(wire714) <<< (~^wire714))}) + $unsigned($signed(((reg720 ?
                  wire706 : reg722) <= $unsigned(wire707)))));
              reg724 <= $unsigned(($signed(reg716[(3'h6):(3'h4)]) ?
                  $signed(reg718[(4'hb):(2'h2)]) : $signed({(wire711 * wire710)})));
            end
          reg725 <= reg716[(1'h1):(1'h0)];
          for (forvar726 = (1'h0); (forvar726 < (2'h3)); forvar726 = (forvar726 + (1'h1)))
            begin
              reg727 = (~(-(+(reg724 > (reg720 ? wire706 : reg717)))));
              reg728 <= (^($signed((^{wire712, reg720})) ^~ reg715));
            end
        end
    end
  assign wire729 = $unsigned(wire707);
  assign wire730 = reg725;
  assign wire731 = (~^reg728[(5'h10):(3'h7)]);
  assign wire732 = (~&$signed($signed(wire706[(1'h0):(1'h0)])));
  assign wire733 = reg728;
  always
    @(posedge clk) begin
      for (forvar734 = (1'h0); (forvar734 < (1'h0)); forvar734 = (forvar734 + (1'h1)))
        begin
          for (forvar735 = (1'h0); (forvar735 < (3'h4)); forvar735 = (forvar735 + (1'h1)))
            begin
              reg736 <= (wire714 << (((((8'hb5) ?
                      wire711 : (8'ha3)) * (wire710 && wire729)) + (^reg728[(4'h8):(3'h7)])) ?
                  wire712[(3'h5):(3'h4)] : (-$signed(wire731))));
              reg737 = $signed(wire712[(3'h4):(1'h0)]);
              reg738 <= wire714;
              reg739 = wire729[(1'h1):(1'h1)];
            end
          reg740 <= $unsigned(((^(+(reg722 ? wire732 : reg719))) ?
              wire713 : {$signed((!reg728)),
                  ($unsigned((8'h9e)) ?
                      (wire731 ? wire706 : wire711) : $unsigned((8'hbd)))}));
          reg741 = wire712;
        end
      reg742 <= (+reg740[(3'h4):(1'h0)]);
      for (forvar743 = (1'h0); (forvar743 < (2'h2)); forvar743 = (forvar743 + (1'h1)))
        begin
          for (forvar744 = (1'h0); (forvar744 < (1'h0)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 <= ($unsigned(wire732[(1'h0):(1'h0)]) * {{$signed({wire729,
                          reg719})},
                  reg741});
              reg746 = (~|(reg722 >> ($signed(forvar735[(4'he):(2'h3)]) & $signed({reg728}))));
              reg747 <= reg740;
              reg748 = {(forvar735[(4'hb):(2'h3)] <= wire713)};
            end
          for (forvar749 = (1'h0); (forvar749 < (1'h1)); forvar749 = (forvar749 + (1'h1)))
            begin
              reg750 <= {$unsigned({((reg724 ? forvar743 : reg737) ?
                          (wire733 & wire732) : forvar734[(2'h2):(2'h2)])})};
              reg751 = ($signed($signed(reg737)) ?
                  (reg742 - $signed(($signed(wire710) ?
                      (reg739 < reg722) : reg737))) : ({reg717,
                          (forvar744[(3'h5):(2'h2)] ?
                              (~^reg728) : $unsigned(reg736))} ?
                      reg737 : wire711));
            end
          reg752 = (reg722 ?
              (~&wire710) : ($unsigned(reg725) ?
                  $signed(((reg725 ? (7'h41) : wire708) >>> {reg741,
                      reg722})) : ((~reg746) ?
                      (reg717 ? (^reg739) : (^~reg736)) : ({reg742} ?
                          (^forvar734) : (~|(8'ha7))))));
          reg753 = $unsigned((!$unsigned(reg738[(4'hb):(3'h4)])));
          if (wire729)
            begin
              reg754 <= ($signed({$unsigned((+wire708))}) ?
                  (-$signed(reg724)) : (($signed(reg740) ?
                      (8'hba) : $unsigned((reg728 ?
                          (8'had) : wire732))) >= $unsigned($signed((~reg736)))));
              reg755 = (~|$unsigned(reg725));
              reg756 <= (wire733[(4'h9):(3'h4)] ?
                  (8'hb0) : (~&($signed(wire731) ?
                      (~|reg717[(5'h12):(3'h7)]) : (^(reg728 | wire712)))));
              reg757 <= $unsigned((({$unsigned(reg722), $unsigned(forvar749)} ?
                  (~^forvar744[(3'h4):(2'h3)]) : {$signed((7'h41))}) & ((8'ha0) ?
                  reg747 : $signed(wire707[(5'h12):(3'h6)]))));
            end
          else
            begin
              reg754 <= $unsigned(reg756[(3'h5):(1'h0)]);
              reg755 = (8'h9e);
            end
        end
      reg758 = (~&$signed($unsigned($unsigned($unsigned(reg725)))));
    end
  assign wire759 = reg740[(4'ha):(3'h4)];
  assign wire760 = $unsigned((wire710[(2'h3):(1'h1)] ^ {reg717[(5'h17):(4'h8)]}));
  assign wire761 = (($signed($signed(wire714)) ?
                       (+(~&$signed(wire707))) : wire733[(4'ha):(2'h2)]) - (wire759[(5'h10):(1'h0)] + $signed((reg725[(3'h7):(2'h3)] & (reg736 ?
                       (8'ha1) : wire729)))));
  always
    @(posedge clk) begin
      reg762 = $unsigned(((((wire730 == wire760) ^~ (reg738 ?
              wire761 : reg728)) ?
          wire707 : wire733) ^~ (~^$unsigned($signed(wire731)))));
      for (forvar763 = (1'h0); (forvar763 < (1'h1)); forvar763 = (forvar763 + (1'h1)))
        begin
          if ((reg719[(1'h0):(1'h0)] >>> $signed($signed((+reg754[(5'h18):(3'h4)])))))
            begin
              reg764 <= (~|$signed({($unsigned((7'h44)) ?
                      (~|wire733) : (wire732 << (7'h40))),
                  reg738}));
              reg765 <= (reg750 ?
                  ((reg725[(5'h14):(4'hf)] ? wire714[(2'h2):(1'h0)] : wire730) ?
                      (reg724 != reg717[(4'hf):(4'hd)]) : reg754[(1'h0):(1'h0)]) : wire706[(2'h2):(2'h2)]);
              reg766 <= (+(7'h40));
              reg767 <= ($signed((reg728[(5'h11):(4'h8)] ?
                      wire761[(2'h3):(1'h0)] : (^wire731))) ?
                  $signed(reg740[(3'h7):(3'h7)]) : {$signed(reg762),
                      (!$unsigned((8'ha8)))});
            end
          else
            begin
              reg764 <= ({reg766[(1'h1):(1'h1)],
                      (~$unsigned(reg766[(1'h1):(1'h0)]))} ?
                  $unsigned({((~wire760) ? $signed(wire761) : (8'hbc)),
                      $unsigned(wire706)}) : reg716[(3'h4):(1'h0)]);
            end
        end
      reg768 = (&reg765);
    end
  assign wire769 = ($unsigned((~|(wire706[(1'h1):(1'h0)] - (reg722 ?
                           (8'hb2) : reg728)))) ?
                       ((^~(!(~wire729))) * wire709) : ($unsigned((^~(~reg754))) ?
                           $signed($signed(reg725[(1'h0):(1'h0)])) : $unsigned(($unsigned(reg757) ?
                               {wire712} : $unsigned(reg725)))));
  always
    @(posedge clk) begin
      reg770 <= (^wire760);
      if ((^~({(~$signed(wire732)), (!(7'h48))} ?
          $signed({(wire706 > wire713),
              (~reg717)}) : (wire730 != $unsigned($signed(reg736))))))
        begin
          reg771 <= ((reg765 != $signed($signed((7'h48)))) > $signed($unsigned((^~(reg750 * wire712)))));
        end
      else
        begin
          for (forvar771 = (1'h0); (forvar771 < (2'h3)); forvar771 = (forvar771 + (1'h1)))
            begin
              reg772 <= reg750;
              reg773 <= $signed({(!reg736[(2'h3):(1'h0)]),
                  ((wire761 ^ (8'hb2)) ? reg716 : reg771)});
              reg774 <= $signed((&wire708));
              reg775 <= reg772[(3'h5):(2'h3)];
            end
        end
      for (forvar776 = (1'h0); (forvar776 < (1'h0)); forvar776 = (forvar776 + (1'h1)))
        begin
          reg777 <= $signed((~&reg774[(4'hc):(4'ha)]));
        end
    end
  always
    @(posedge clk) begin
      reg778 <= (~|(~wire769));
    end
  always
    @(posedge clk) begin
      for (forvar779 = (1'h0); (forvar779 < (1'h0)); forvar779 = (forvar779 + (1'h1)))
        begin
          reg780 = $signed(({reg745,
              $signed($unsigned(wire712))} < $unsigned($unsigned((forvar779 >> reg771)))));
          reg781 = reg724[(3'h6):(1'h0)];
        end
      reg782 = (^~(|(!reg766)));
      if ({wire760[(3'h7):(1'h1)], (&(~reg765))})
        begin
          for (forvar783 = (1'h0); (forvar783 < (2'h3)); forvar783 = (forvar783 + (1'h1)))
            begin
              reg784 <= wire710[(2'h2):(2'h2)];
              reg785 = $unsigned((|((8'hb6) > $unsigned($unsigned(reg766)))));
              reg786 = $signed(reg722);
              reg787 = {reg738[(3'h6):(1'h1)], $unsigned(wire769)};
            end
          reg788 = $signed(reg757);
          if (wire712)
            begin
              reg789 = reg777[(2'h3):(1'h0)];
              reg790 = reg770;
            end
          else
            begin
              reg789 = (forvar783[(4'h9):(2'h3)] ?
                  (8'ha3) : ((wire761[(3'h5):(1'h1)] ? reg767 : (8'h9f)) ?
                      (~^reg770[(4'ha):(3'h4)]) : (((wire730 - reg736) >>> $unsigned(wire731)) && $unsigned(((7'h49) ?
                          reg717 : reg736)))));
            end
        end
      else
        begin
          for (forvar783 = (1'h0); (forvar783 < (2'h3)); forvar783 = (forvar783 + (1'h1)))
            begin
              reg784 <= {$signed($unsigned((8'ha4))),
                  (|(reg724 || $unsigned((reg767 ? reg773 : wire713))))};
              reg791 <= (~^(reg740 ?
                  (~reg725) : ({(reg764 < wire713)} ?
                      wire707[(5'h17):(2'h3)] : ($unsigned(wire706) ?
                          {reg764} : (wire710 >>> reg784)))));
              reg792 <= reg773[(4'hc):(3'h4)];
            end
        end
      for (forvar793 = (1'h0); (forvar793 < (3'h4)); forvar793 = (forvar793 + (1'h1)))
        begin
          reg794 = (&reg777);
          if (wire709)
            begin
              reg795 <= reg754;
            end
          else
            begin
              reg795 <= ((8'hba) >>> ((((wire759 ^~ reg736) ^~ $signed(wire714)) > ($signed((8'ha8)) ?
                      (8'hb4) : $unsigned(wire706))) ?
                  reg754 : reg772[(3'h4):(1'h1)]));
              reg796 <= wire729;
            end
        end
    end
  assign wire797 = (-wire713);
  assign wire798 = $unsigned(wire759[(4'he):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module446  (y, clk, wire450, wire449, wire448, wire447);
  output wire [(32'hd11):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h16):(1'h0)] wire450;
  input wire signed [(4'hf):(1'h0)] wire449;
  input wire [(4'hb):(1'h0)] wire448;
  input wire signed [(5'h12):(1'h0)] wire447;
  wire [(3'h5):(1'h0)] wire659;
  wire signed [(4'hf):(1'h0)] wire658;
  wire signed [(4'h8):(1'h0)] wire646;
  wire signed [(4'hf):(1'h0)] wire645;
  wire [(3'h5):(1'h0)] wire643;
  wire signed [(5'h12):(1'h0)] wire618;
  wire signed [(5'h18):(1'h0)] wire617;
  wire [(4'ha):(1'h0)] wire616;
  wire signed [(4'he):(1'h0)] wire587;
  wire [(5'h11):(1'h0)] wire564;
  wire signed [(3'h5):(1'h0)] wire563;
  wire [(3'h7):(1'h0)] wire562;
  wire [(2'h2):(1'h0)] wire561;
  wire signed [(5'h14):(1'h0)] wire560;
  reg [(3'h5):(1'h0)] reg683 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg681 = (1'h0);
  reg [(3'h4):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg691 = (1'h0);
  reg [(2'h3):(1'h0)] reg690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg685 = (1'h0);
  reg [(3'h7):(1'h0)] reg684 = (1'h0);
  reg [(5'h17):(1'h0)] reg680 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg678 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg674 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg673 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg670 = (1'h0);
  reg [(4'h9):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg657 = (1'h0);
  reg [(4'hb):(1'h0)] reg653 = (1'h0);
  reg [(5'h12):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg648 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg644 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg641 = (1'h0);
  reg [(5'h17):(1'h0)] reg639 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg634 = (1'h0);
  reg [(2'h2):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg630 = (1'h0);
  reg signed [(4'he):(1'h0)] reg625 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg624 = (1'h0);
  reg [(5'h13):(1'h0)] reg623 = (1'h0);
  reg [(4'he):(1'h0)] reg620 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg619 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg615 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg613 = (1'h0);
  reg [(3'h7):(1'h0)] reg612 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg611 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg609 = (1'h0);
  reg [(2'h3):(1'h0)] reg607 = (1'h0);
  reg [(4'h8):(1'h0)] reg606 = (1'h0);
  reg [(4'hc):(1'h0)] reg604 = (1'h0);
  reg [(5'h17):(1'h0)] reg603 = (1'h0);
  reg [(3'h4):(1'h0)] reg601 = (1'h0);
  reg [(5'h16):(1'h0)] reg588 = (1'h0);
  reg [(2'h3):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg594 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg592 = (1'h0);
  reg [(4'hc):(1'h0)] reg591 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg590 = (1'h0);
  reg [(4'hb):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg583 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg582 = (1'h0);
  reg [(4'hf):(1'h0)] reg576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg572 = (1'h0);
  reg [(5'h16):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg569 = (1'h0);
  reg [(5'h18):(1'h0)] reg567 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg565 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg556 = (1'h0);
  reg [(5'h18):(1'h0)] reg552 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg550 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg549 = (1'h0);
  reg [(5'h12):(1'h0)] reg547 = (1'h0);
  reg signed [(4'he):(1'h0)] reg546 = (1'h0);
  reg [(4'hc):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg542 = (1'h0);
  reg [(4'h8):(1'h0)] reg541 = (1'h0);
  reg [(4'hd):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg536 = (1'h0);
  reg [(4'h8):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg527 = (1'h0);
  reg [(5'h18):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg525 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg524 = (1'h0);
  reg [(4'he):(1'h0)] reg520 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg518 = (1'h0);
  reg signed [(4'he):(1'h0)] reg513 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg510 = (1'h0);
  reg [(4'hb):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg506 = (1'h0);
  reg [(2'h3):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg504 = (1'h0);
  reg [(4'h8):(1'h0)] reg503 = (1'h0);
  reg [(5'h13):(1'h0)] reg502 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg500 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg494 = (1'h0);
  reg [(5'h11):(1'h0)] reg492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg489 = (1'h0);
  reg [(4'h9):(1'h0)] reg488 = (1'h0);
  reg [(5'h10):(1'h0)] reg486 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg483 = (1'h0);
  reg [(2'h2):(1'h0)] reg480 = (1'h0);
  reg [(5'h18):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg477 = (1'h0);
  reg [(5'h10):(1'h0)] reg473 = (1'h0);
  reg [(4'hc):(1'h0)] reg472 = (1'h0);
  reg [(5'h10):(1'h0)] reg467 = (1'h0);
  reg [(4'h8):(1'h0)] reg466 = (1'h0);
  reg [(4'hb):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg461 = (1'h0);
  reg [(3'h4):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg457 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg455 = (1'h0);
  reg [(4'hd):(1'h0)] reg452 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg692 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar679 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar675 = (1'h0);
  reg [(3'h4):(1'h0)] forvar692 = (1'h0);
  reg [(5'h10):(1'h0)] reg689 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar683 = (1'h0);
  reg [(5'h17):(1'h0)] reg682 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar681 = (1'h0);
  reg [(4'h8):(1'h0)] reg679 = (1'h0);
  reg [(4'hb):(1'h0)] reg677 = (1'h0);
  reg [(3'h6):(1'h0)] reg676 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg675 = (1'h0);
  reg [(4'hc):(1'h0)] reg672 = (1'h0);
  reg [(4'hd):(1'h0)] forvar671 = (1'h0);
  reg [(5'h12):(1'h0)] reg669 = (1'h0);
  reg [(5'h14):(1'h0)] forvar668 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg664 = (1'h0);
  reg [(5'h17):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar662 = (1'h0);
  reg [(3'h7):(1'h0)] forvar661 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg660 = (1'h0);
  reg [(4'h8):(1'h0)] reg656 = (1'h0);
  reg [(5'h10):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg654 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar652 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg650 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar649 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg647 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg636 = (1'h0);
  reg [(5'h14):(1'h0)] forvar635 = (1'h0);
  reg [(5'h16):(1'h0)] forvar633 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg629 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar627 = (1'h0);
  reg [(5'h18):(1'h0)] reg626 = (1'h0);
  reg [(5'h16):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg621 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg614 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar608 = (1'h0);
  reg [(3'h5):(1'h0)] forvar604 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg602 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg599 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg598 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar596 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg595 = (1'h0);
  reg [(4'h8):(1'h0)] reg593 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg589 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar588 = (1'h0);
  reg [(4'he):(1'h0)] reg585 = (1'h0);
  reg [(2'h2):(1'h0)] reg584 = (1'h0);
  reg [(5'h12):(1'h0)] reg581 = (1'h0);
  reg [(5'h16):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar579 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg578 = (1'h0);
  reg [(4'hc):(1'h0)] reg577 = (1'h0);
  reg [(3'h4):(1'h0)] reg575 = (1'h0);
  reg [(5'h18):(1'h0)] reg574 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar572 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg573 = (1'h0);
  reg [(4'hd):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg566 = (1'h0);
  reg [(4'he):(1'h0)] reg555 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg554 = (1'h0);
  reg [(4'h9):(1'h0)] reg553 = (1'h0);
  reg [(4'h9):(1'h0)] forvar551 = (1'h0);
  reg [(5'h12):(1'h0)] reg548 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg545 = (1'h0);
  reg [(4'he):(1'h0)] reg544 = (1'h0);
  reg [(5'h17):(1'h0)] forvar540 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg539 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg537 = (1'h0);
  reg [(3'h7):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar534 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar533 = (1'h0);
  reg [(4'hc):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg523 = (1'h0);
  reg [(4'hb):(1'h0)] reg522 = (1'h0);
  reg [(5'h16):(1'h0)] forvar521 = (1'h0);
  reg [(4'h8):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar517 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg515 = (1'h0);
  reg [(4'he):(1'h0)] forvar514 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg512 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg511 = (1'h0);
  reg [(4'hd):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg501 = (1'h0);
  reg [(3'h5):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar498 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg497 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg496 = (1'h0);
  reg [(3'h5):(1'h0)] reg495 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar493 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg491 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg490 = (1'h0);
  reg [(5'h10):(1'h0)] reg487 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg484 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar478 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg476 = (1'h0);
  reg [(5'h11):(1'h0)] forvar475 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg471 = (1'h0);
  reg [(5'h15):(1'h0)] reg470 = (1'h0);
  reg [(5'h17):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg468 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg465 = (1'h0);
  reg [(3'h4):(1'h0)] forvar463 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg460 = (1'h0);
  reg signed [(4'he):(1'h0)] reg453 = (1'h0);
  reg [(4'h9):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg454 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar453 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg451 = (1'h0);
  assign y = {wire659,
                 wire658,
                 wire646,
                 wire645,
                 wire643,
                 wire618,
                 wire617,
                 wire616,
                 wire587,
                 wire564,
                 wire563,
                 wire562,
                 wire561,
                 wire560,
                 reg683,
                 reg681,
                 reg693,
                 reg691,
                 reg690,
                 reg688,
                 reg685,
                 reg684,
                 reg680,
                 reg678,
                 reg674,
                 reg673,
                 reg670,
                 reg667,
                 reg666,
                 reg665,
                 reg657,
                 reg653,
                 reg651,
                 reg648,
                 reg644,
                 reg641,
                 reg639,
                 reg638,
                 reg637,
                 reg634,
                 reg631,
                 reg630,
                 reg625,
                 reg624,
                 reg623,
                 reg620,
                 reg619,
                 reg615,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg607,
                 reg606,
                 reg604,
                 reg603,
                 reg601,
                 reg588,
                 reg597,
                 reg594,
                 reg592,
                 reg591,
                 reg590,
                 reg586,
                 reg583,
                 reg582,
                 reg576,
                 reg572,
                 reg571,
                 reg569,
                 reg567,
                 reg565,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg552,
                 reg550,
                 reg549,
                 reg547,
                 reg546,
                 reg543,
                 reg542,
                 reg541,
                 reg538,
                 reg536,
                 reg532,
                 reg531,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg520,
                 reg518,
                 reg513,
                 reg510,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg500,
                 reg494,
                 reg492,
                 reg489,
                 reg488,
                 reg486,
                 reg483,
                 reg480,
                 reg479,
                 reg477,
                 reg473,
                 reg472,
                 reg467,
                 reg466,
                 reg464,
                 reg461,
                 reg459,
                 reg457,
                 reg456,
                 reg455,
                 reg452,
                 reg692,
                 forvar679,
                 forvar675,
                 forvar692,
                 reg689,
                 reg687,
                 reg686,
                 forvar683,
                 reg682,
                 forvar681,
                 reg679,
                 reg677,
                 reg676,
                 reg675,
                 reg672,
                 forvar671,
                 reg669,
                 forvar668,
                 reg664,
                 reg663,
                 forvar662,
                 forvar661,
                 reg660,
                 reg656,
                 reg655,
                 reg654,
                 forvar652,
                 reg650,
                 forvar649,
                 reg647,
                 reg642,
                 reg640,
                 reg636,
                 forvar635,
                 forvar633,
                 reg632,
                 reg629,
                 reg628,
                 forvar627,
                 reg626,
                 reg622,
                 reg621,
                 reg614,
                 forvar608,
                 forvar604,
                 reg605,
                 reg602,
                 reg600,
                 reg599,
                 reg598,
                 forvar596,
                 reg595,
                 reg593,
                 reg589,
                 forvar588,
                 reg585,
                 reg584,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg577,
                 reg575,
                 reg574,
                 forvar572,
                 reg573,
                 reg570,
                 reg568,
                 reg566,
                 reg555,
                 reg554,
                 reg553,
                 forvar551,
                 reg548,
                 reg545,
                 reg544,
                 forvar540,
                 reg539,
                 reg537,
                 reg535,
                 forvar534,
                 forvar533,
                 reg530,
                 reg529,
                 reg528,
                 reg523,
                 reg522,
                 forvar521,
                 reg519,
                 forvar517,
                 reg516,
                 reg515,
                 forvar514,
                 reg512,
                 reg511,
                 reg509,
                 reg508,
                 reg501,
                 reg499,
                 forvar498,
                 reg497,
                 reg496,
                 reg495,
                 forvar493,
                 reg491,
                 reg490,
                 reg487,
                 reg485,
                 reg484,
                 reg482,
                 reg481,
                 forvar478,
                 reg476,
                 forvar475,
                 reg474,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg465,
                 forvar463,
                 reg462,
                 reg460,
                 reg453,
                 reg458,
                 reg454,
                 forvar453,
                 reg451,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($unsigned({$unsigned($signed((8'haa))),
              (~&(wire447 ? wire450 : wire448))}) ?
          $unsigned((^~(wire448 ?
              ((8'hbd) ?
                  wire448 : wire447) : wire450))) : {(|$unsigned({wire449,
                  wire447}))}))
        begin
          reg451 = wire448[(2'h3):(1'h1)];
          reg452 <= {$signed(((~^wire449[(4'hf):(1'h1)]) & {$unsigned((7'h45)),
                  $unsigned(wire450)})),
              ($unsigned((wire449 ?
                  $signed(wire449) : (wire448 ^ wire450))) ~^ $unsigned(wire448[(2'h2):(1'h1)]))};
          for (forvar453 = (1'h0); (forvar453 < (3'h4)); forvar453 = (forvar453 + (1'h1)))
            begin
              reg454 = (^(~&(wire448[(4'hb):(3'h4)] ?
                  wire448[(4'hb):(3'h5)] : $unsigned($unsigned(reg452)))));
            end
          if (wire447[(1'h1):(1'h0)])
            begin
              reg455 <= $unsigned({$unsigned((~|(~|reg452))), wire449});
              reg456 <= wire449[(2'h3):(1'h1)];
              reg457 <= (wire447 << $signed((~|($signed(reg452) | wire447[(1'h0):(1'h0)]))));
              reg458 = $signed((reg452 <= {((|forvar453) ?
                      $signed((7'h42)) : $unsigned((8'ha3))),
                  {(8'haf)}}));
            end
          else
            begin
              reg455 <= {reg454,
                  (~|$signed((reg458[(3'h7):(2'h2)] ^ $unsigned(wire450))))};
              reg456 <= (($unsigned($signed((forvar453 >= wire449))) ?
                  (~^wire447) : $unsigned((~|(8'h9c)))) <= {(reg457 & $unsigned((+reg457))),
                  {$signed((wire447 ? wire447 : reg451))}});
              reg457 <= wire447[(3'h4):(3'h4)];
              reg459 <= forvar453;
            end
        end
      else
        begin
          if (($unsigned(reg455) || ($unsigned((~&(wire450 == wire450))) ?
              $unsigned(reg451[(3'h5):(1'h1)]) : (^reg454))))
            begin
              reg451 = reg452[(4'h8):(3'h5)];
              reg453 = (+{(&$signed(wire448)),
                  {wire450,
                      ((reg458 * reg451) ?
                          $signed(wire447) : (reg458 ? reg454 : reg458))}});
              reg455 <= $unsigned(($signed(reg453[(4'hc):(3'h4)]) >> (7'h45)));
              reg458 = ($signed(forvar453[(1'h0):(1'h0)]) - $signed(($signed($unsigned(reg456)) && ({reg459} ?
                  (reg458 ? wire447 : wire449) : reg452))));
            end
          else
            begin
              reg452 <= {(((^(wire450 == reg455)) ?
                      $signed($signed(reg454)) : (^$signed(wire449))) >>> (~|wire447[(3'h7):(1'h1)]))};
              reg453 = ((((7'h4a) ?
                          $signed((wire449 == reg453)) : reg458[(3'h6):(1'h0)]) ?
                      $signed({$unsigned(reg459)}) : ($unsigned($signed(reg452)) ?
                          (^~(!(8'hba))) : $unsigned(reg456))) ?
                  (((-(reg459 ? reg459 : reg458)) ~^ ((8'haa) ?
                      (reg453 <<< reg455) : {(8'hbf)})) - $signed((wire447 ?
                      (-wire449) : reg455))) : {(reg459 != (&{forvar453})),
                      wire450[(4'hf):(4'h8)]});
            end
          if (wire448)
            begin
              reg459 <= (wire449 ^~ (wire450 * $unsigned(((|wire449) == $signed(reg456)))));
              reg460 = $signed(reg453[(4'ha):(3'h7)]);
            end
          else
            begin
              reg460 = (wire449 ?
                  (((reg454 ?
                      wire447 : $signed((8'ha9))) | ((reg460 ^ (8'hb8)) ~^ (wire449 != (7'h48)))) ^~ ((|$signed(reg452)) ?
                      $signed($signed(reg452)) : (|$unsigned(reg451)))) : reg452);
            end
          reg461 <= {wire449, $signed({{{reg459}}})};
          reg462 = {wire447[(4'he):(3'h4)]};
        end
      for (forvar463 = (1'h0); (forvar463 < (1'h1)); forvar463 = (forvar463 + (1'h1)))
        begin
          reg464 <= (reg452 ? reg452 : reg462);
          if ($unsigned($signed((reg460 ? reg453 : reg462[(3'h6):(3'h6)]))))
            begin
              reg465 = $signed($unsigned($signed($unsigned((wire449 ?
                  (8'hb9) : (8'ha8))))));
              reg466 <= (!(wire449[(4'hf):(2'h3)] ? reg453 : reg454));
            end
          else
            begin
              reg466 <= reg466[(1'h1):(1'h0)];
            end
          if ({(forvar463 & {((~&reg457) <= reg460[(5'h17):(4'hd)])})})
            begin
              reg467 <= (&(reg454[(1'h1):(1'h1)] ?
                  $unsigned($signed(forvar453[(1'h0):(1'h0)])) : {$signed($unsigned((8'ha9))),
                      ((reg466 ? reg461 : reg462) != (wire447 ?
                          (8'ha7) : forvar463))}));
              reg468 = (^wire450[(4'he):(4'ha)]);
              reg469 = ((reg455[(3'h4):(1'h0)] ?
                      $unsigned($signed(reg462[(1'h1):(1'h0)])) : wire449[(4'hc):(1'h1)]) ?
                  $unsigned({(~(~|(8'ha7))),
                      {(reg468 && (8'haf)),
                          $signed(reg455)}}) : ((|$signed($unsigned(reg461))) ?
                      (wire448[(3'h5):(1'h1)] * (~^(~^reg465))) : ($unsigned(forvar463) ?
                          reg458 : $unsigned(reg467))));
              reg470 = $signed((8'hbe));
              reg471 = (reg465 ?
                  (~^(((reg452 || reg455) ^~ (-(8'h9f))) && (reg467[(1'h0):(1'h0)] <= (reg461 ?
                      (8'had) : reg462)))) : {({(reg452 && forvar463)} <= {reg470})});
            end
          else
            begin
              reg468 = $signed($signed(reg452[(4'h9):(3'h5)]));
              reg472 <= $signed(reg460[(5'h16):(4'h8)]);
              reg473 <= reg453[(3'h4):(1'h0)];
              reg474 = (&$unsigned((+{reg459[(2'h3):(2'h3)],
                  ((7'h42) <= wire450)})));
            end
          for (forvar475 = (1'h0); (forvar475 < (1'h0)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 = $unsigned(reg459);
              reg477 <= {(((8'hae) >>> $signed($unsigned(forvar453))) + reg451)};
            end
          for (forvar478 = (1'h0); (forvar478 < (2'h3)); forvar478 = (forvar478 + (1'h1)))
            begin
              reg479 <= (|(forvar475[(3'h7):(3'h5)] < {reg457,
                  {(reg472 >>> wire447)}}));
              reg480 <= (~|reg459);
              reg481 = reg480[(2'h2):(2'h2)];
              reg482 = $unsigned($unsigned($unsigned(wire449)));
              reg483 <= (~|($unsigned((^~(reg471 > reg481))) ?
                  (^reg464[(1'h1):(1'h0)]) : $unsigned($signed(reg454))));
            end
        end
      reg484 = reg465;
      reg485 = {reg452[(1'h0):(1'h0)], wire447};
      if (($unsigned(($unsigned($signed(reg477)) ?
          (forvar453 <<< $unsigned(reg453)) : ((~wire447) <<< (+(8'hbb))))) >>> {(+($unsigned(reg467) ?
              $unsigned(wire448) : $signed((8'h9f)))),
          (~&{(!reg485), $signed((8'hae))})}))
        begin
          reg486 <= reg456;
          reg487 = $unsigned($unsigned((~forvar463)));
          if (reg471)
            begin
              reg488 <= reg461[(1'h0):(1'h0)];
              reg489 <= $signed({(reg455 ?
                      ((forvar478 && (7'h43)) ?
                          reg471 : (8'h9e)) : reg466[(1'h0):(1'h0)])});
              reg490 = (8'ha3);
              reg491 = $unsigned(wire450[(2'h3):(1'h1)]);
            end
          else
            begin
              reg488 <= {(forvar475[(3'h6):(1'h1)] || (!((reg476 ?
                          reg481 : reg482) ?
                      $unsigned(reg477) : ((8'hb4) - reg467)))),
                  $unsigned(reg459)};
              reg490 = {{reg468[(4'hc):(2'h3)], wire447},
                  (!(~|reg473[(2'h2):(1'h0)]))};
            end
          reg492 <= (8'hb7);
          for (forvar493 = (1'h0); (forvar493 < (2'h2)); forvar493 = (forvar493 + (1'h1)))
            begin
              reg494 <= reg476[(2'h3):(2'h2)];
              reg495 = (~(($signed($signed(reg454)) || reg481) ?
                  $unsigned(($unsigned(reg455) * $unsigned(forvar478))) : reg471[(3'h5):(3'h5)]));
              reg496 = (reg454[(3'h6):(1'h1)] ?
                  $signed($signed((reg495 ?
                      reg459[(2'h2):(1'h1)] : (reg452 ^ reg489)))) : $unsigned($signed((reg480 ?
                      forvar453[(1'h1):(1'h0)] : {reg451, (8'ha9)}))));
              reg497 = ((!(forvar463[(2'h2):(2'h2)] < (|$unsigned(reg458)))) ?
                  (^(reg479 > reg468[(4'h9):(1'h0)])) : {($unsigned($unsigned(reg471)) << ((reg489 ?
                              reg471 : forvar478) ?
                          $signed(reg496) : $signed(reg459))),
                      ({reg473[(4'h8):(3'h7)], wire449[(3'h5):(2'h2)]} ?
                          ({reg483, reg459} ?
                              (|reg453) : (reg451 ?
                                  reg467 : reg466)) : reg492)});
            end
        end
      else
        begin
          reg487 = (~^reg469[(5'h13):(3'h5)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar498 = (1'h0); (forvar498 < (3'h4)); forvar498 = (forvar498 + (1'h1)))
        begin
          if (reg452)
            begin
              reg499 = $signed({{($unsigned(reg494) ?
                          (wire448 == wire449) : $signed(reg477))},
                  (-((8'hac) ?
                      (forvar498 ?
                          (7'h46) : reg480) : wire448[(3'h4):(1'h0)]))});
              reg500 <= reg480;
              reg501 = (8'hb9);
            end
          else
            begin
              reg499 = reg494;
              reg501 = wire449;
              reg502 <= reg473;
              reg503 <= (-(8'h9f));
            end
          if (forvar498[(4'hf):(1'h0)])
            begin
              reg504 <= wire448;
              reg505 <= (!((&forvar498) << (~^$unsigned((~^reg466)))));
              reg506 <= ($signed(reg457[(1'h0):(1'h0)]) ?
                  (!$unsigned($unsigned(forvar498[(3'h6):(3'h6)]))) : reg489);
              reg507 <= (reg499[(2'h2):(1'h0)] < wire449);
              reg508 = (((|reg459[(1'h0):(1'h0)]) ?
                      $unsigned($unsigned((&reg507))) : (({reg503} << $unsigned(reg500)) >>> ((reg494 * reg480) ?
                          reg464 : reg505[(2'h3):(1'h1)]))) ?
                  (reg452 >>> ($unsigned((reg466 ? reg466 : reg500)) ?
                      {{reg477, reg467},
                          (reg452 ?
                              (8'ha0) : forvar498)} : wire450)) : $signed($unsigned({reg452[(2'h2):(1'h0)],
                      (8'hbe)})));
            end
          else
            begin
              reg508 = wire449[(3'h7):(3'h4)];
              reg509 = reg472[(2'h2):(2'h2)];
              reg510 <= (8'ha5);
              reg511 = ((($signed((~^reg503)) ?
                      $unsigned(reg479[(3'h5):(2'h3)]) : ($unsigned((8'ha8)) < (reg483 ?
                          (8'hbc) : wire449))) ?
                  {(7'h46),
                      ({reg500, reg479} ?
                          reg503 : (wire450 ?
                              reg472 : wire448))} : (^(wire450 && $unsigned((8'h9f))))) >>> $signed($unsigned(($unsigned(reg479) | (reg466 ?
                  reg492 : reg480)))));
            end
          reg512 = (reg502 <= (reg508[(2'h2):(1'h0)] | wire447[(5'h12):(4'hc)]));
          reg513 <= $signed(reg489[(1'h0):(1'h0)]);
        end
      for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
        begin
          reg515 = (+reg509[(4'h9):(3'h5)]);
          reg516 = {($signed($signed({reg508, reg472})) ?
                  (wire448[(1'h1):(1'h0)] ?
                      reg479 : reg455) : reg472[(4'ha):(3'h5)]),
              ($signed((~&forvar498[(5'h15):(4'hd)])) + (reg467[(2'h3):(2'h3)] << $signed(reg503[(1'h1):(1'h0)])))};
          for (forvar517 = (1'h0); (forvar517 < (1'h1)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 <= (reg477 ?
                  $signed(reg511) : $signed($signed($signed(reg516))));
              reg519 = reg510;
              reg520 <= $signed(($unsigned(reg505) && $signed($signed($unsigned(reg486)))));
            end
          for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 = ($unsigned(((^~reg510) ?
                  $unsigned(forvar498) : reg486[(3'h7):(2'h3)])) == ((reg516 * (^~{reg480})) ?
                  forvar514[(2'h3):(2'h3)] : reg518));
              reg523 = (8'ha4);
              reg524 <= ({$signed(($unsigned((7'h41)) & reg486[(1'h1):(1'h0)]))} * {$unsigned($signed((reg515 - wire448)))});
              reg525 <= $unsigned(forvar521[(5'h11):(1'h0)]);
            end
        end
      if ((reg507 ? reg513[(1'h1):(1'h0)] : reg501[(5'h12):(2'h3)]))
        begin
          reg526 <= (reg511[(1'h0):(1'h0)] & $unsigned($unsigned(({reg486} + $unsigned(reg473)))));
          reg527 <= reg509;
          reg528 = $signed(reg509);
        end
      else
        begin
          reg526 <= $signed(reg492[(3'h7):(3'h4)]);
          reg527 <= reg526;
          reg528 = ((^~$unsigned(reg492)) || {$signed(forvar517)});
          reg529 = (~&reg473[(1'h0):(1'h0)]);
          if (($signed(((^~((8'hb6) - reg452)) ?
                  reg499[(2'h2):(2'h2)] : $unsigned((reg516 ^~ reg494)))) ?
              $signed((^$signed((-reg492)))) : reg524[(1'h0):(1'h0)]))
            begin
              reg530 = ((!{(reg528[(4'ha):(2'h2)] ?
                          reg518[(1'h0):(1'h0)] : {reg516, reg502})}) ?
                  $unsigned(reg528[(2'h3):(1'h1)]) : ({$unsigned((~reg519)),
                      ({reg457} * {reg459, reg452})} <<< $unsigned({reg504})));
              reg531 <= reg526;
            end
          else
            begin
              reg530 = (($signed((reg528 >>> $unsigned(reg483))) < (reg520[(3'h7):(1'h1)] <<< reg525[(3'h6):(2'h3)])) || $signed(reg477[(1'h0):(1'h0)]));
              reg531 <= $unsigned(reg509);
              reg532 <= $unsigned((~&(~$unsigned(((8'hba) - reg528)))));
            end
        end
      for (forvar533 = (1'h0); (forvar533 < (2'h3)); forvar533 = (forvar533 + (1'h1)))
        begin
          for (forvar534 = (1'h0); (forvar534 < (3'h4)); forvar534 = (forvar534 + (1'h1)))
            begin
              reg535 = wire448;
              reg536 <= {(!(({reg527, (8'ha6)} ?
                      {(8'hb6)} : reg526) + ((|reg503) ? reg505 : (~|reg520)))),
                  (($signed(reg525) ?
                          (^~(~|reg486)) : (reg459[(1'h1):(1'h0)] != $unsigned(wire447))) ?
                      $unsigned((~^reg535[(3'h5):(3'h4)])) : reg509[(2'h2):(1'h1)])};
            end
          reg537 = reg520;
          if ($signed($unsigned((~^$signed((reg506 <= wire449))))))
            begin
              reg538 <= forvar498[(4'hc):(3'h7)];
            end
          else
            begin
              reg539 = reg527;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar540 = (1'h0); (forvar540 < (3'h4)); forvar540 = (forvar540 + (1'h1)))
        begin
          if ($unsigned($unsigned((reg489[(3'h4):(1'h0)] - reg464))))
            begin
              reg541 <= $signed({($unsigned(reg467[(4'hc):(1'h1)]) | $unsigned((~|wire448))),
                  $unsigned(((wire449 * forvar540) ?
                      reg513[(2'h2):(2'h2)] : (reg477 && reg513)))});
            end
          else
            begin
              reg541 <= $unsigned($unsigned(($signed(reg503[(4'h8):(3'h5)]) < (reg456[(2'h3):(2'h2)] >> $signed(reg510)))));
            end
          if ({{reg480}})
            begin
              reg542 <= ($unsigned(reg518[(1'h1):(1'h1)]) == reg492);
              reg543 <= (~|$signed($signed(reg526[(2'h2):(1'h1)])));
            end
          else
            begin
              reg542 <= reg541;
              reg544 = wire448;
              reg545 = $unsigned($unsigned(($signed({reg518}) & $unsigned((reg506 | reg455)))));
              reg546 <= ({({((8'ha4) >> reg507), (wire450 < reg506)} ?
                      $unsigned((reg543 ? reg504 : reg486)) : reg488),
                  (~((reg489 ? wire447 : reg507) > (reg500 ?
                      reg503 : reg507)))} == reg544[(3'h6):(2'h3)]);
            end
          if ($unsigned($unsigned($unsigned({$signed(reg466),
              (reg527 * reg464)}))))
            begin
              reg547 <= ((8'hb6) ?
                  (reg502[(2'h2):(2'h2)] ?
                      $signed(($signed(reg518) ?
                          reg507 : (reg480 > reg459))) : reg456) : reg502);
              reg548 = ((^$signed(reg480[(2'h2):(2'h2)])) ?
                  (-(({reg513} ?
                      (reg472 && reg494) : $unsigned(reg527)) && (reg542 | reg483[(2'h3):(1'h1)]))) : ({(~^(wire450 >>> reg544))} ^~ {((reg513 ~^ reg480) + $signed(reg536))}));
            end
          else
            begin
              reg547 <= reg541;
              reg548 = ($signed((reg548[(5'h12):(4'h8)] ?
                  (reg459 + (~&(8'hb5))) : {$unsigned((8'ha4))})) ^ ({$signed(wire448)} >= (reg488 <= reg483[(4'he):(4'he)])));
              reg549 <= (+reg503[(1'h0):(1'h0)]);
            end
          reg550 <= $signed($signed({$signed(reg467[(3'h6):(3'h6)]),
              $signed((7'h40))}));
        end
      for (forvar551 = (1'h0); (forvar551 < (3'h4)); forvar551 = (forvar551 + (1'h1)))
        begin
          if (reg542)
            begin
              reg552 <= (-reg506);
              reg553 = reg492;
              reg554 = $unsigned($unsigned($unsigned(reg455)));
              reg555 = ({reg545, ((~|(reg531 + reg452)) & $unsigned(reg506))} ?
                  reg548 : (~(-{$unsigned(reg554)})));
            end
          else
            begin
              reg552 <= ((((8'ha1) <<< reg452) ?
                  $signed(reg546[(3'h4):(1'h0)]) : reg543[(3'h4):(3'h4)]) - reg531[(1'h1):(1'h1)]);
              reg553 = reg492[(4'ha):(1'h1)];
              reg556 <= (($unsigned($unsigned($unsigned((8'had)))) ?
                  $signed((^~reg549)) : ({{reg548}, $unsigned(reg527)} ?
                      (~|reg459) : ((reg544 ? reg520 : reg504) ?
                          (reg548 <= reg507) : reg518))) == {$unsigned(reg553)});
              reg557 <= $signed((~^$unsigned($unsigned(reg547))));
              reg558 <= reg492;
            end
          reg559 <= (((8'ha3) < (8'ha9)) ? reg520 : reg556);
        end
    end
  assign wire560 = $unsigned(reg550[(2'h2):(2'h2)]);
  assign wire561 = $unsigned(reg505[(1'h1):(1'h0)]);
  assign wire562 = reg547[(2'h2):(1'h1)];
  assign wire563 = {$signed({$signed({reg543, reg513}), (^~reg559)})};
  assign wire564 = $signed(reg472[(4'hc):(4'hc)]);
  always
    @(posedge clk) begin
      if ((8'hb9))
        begin
          if ((((8'hb1) ?
              reg461 : $signed((~{reg546}))) << reg502[(4'hd):(1'h0)]))
            begin
              reg565 <= $unsigned(reg486[(4'he):(3'h5)]);
            end
          else
            begin
              reg565 <= reg556[(5'h10):(4'h9)];
              reg566 = wire447;
              reg567 <= (reg520 ? reg480[(1'h1):(1'h1)] : (^reg525));
              reg568 = {(reg542[(1'h0):(1'h0)] > (~{{wire448}, (~^reg527)})),
                  $unsigned((wire560 ? reg558 : $signed((reg532 >> reg455))))};
            end
          reg569 <= $unsigned((8'h9f));
        end
      else
        begin
          if (wire561)
            begin
              reg565 <= (~|reg467);
              reg567 <= reg473[(2'h3):(2'h2)];
              reg569 <= reg502;
              reg570 = ({reg479} ?
                  wire449[(3'h4):(1'h0)] : reg489[(1'h0):(1'h0)]);
            end
          else
            begin
              reg566 = (8'hb6);
            end
        end
      reg571 <= wire561;
      if (wire560[(4'hd):(1'h1)])
        begin
          reg572 <= $unsigned((($unsigned((~reg500)) ?
              reg459 : reg502[(4'h9):(1'h0)]) & {$signed(((8'ha6) * reg550))}));
          reg573 = $signed((($signed({(8'ha0), wire560}) ?
                  reg566[(4'h9):(1'h1)] : {$signed(reg452), (~^reg543)}) ?
              $unsigned(((reg558 ?
                  (8'haf) : reg494) >> (reg572 || reg505))) : {$signed($unsigned(wire563)),
                  $unsigned($unsigned(reg538))}));
        end
      else
        begin
          for (forvar572 = (1'h0); (forvar572 < (1'h1)); forvar572 = (forvar572 + (1'h1)))
            begin
              reg573 = reg506[(4'hb):(3'h4)];
            end
          if ($signed((!$signed(reg559[(2'h2):(2'h2)]))))
            begin
              reg574 = (((reg557[(3'h5):(1'h1)] ^~ ((reg507 * reg541) ?
                          (reg467 ?
                              reg538 : (8'haf)) : reg558[(3'h7):(3'h4)])) ?
                      {(8'ha6),
                          (reg486[(4'hf):(3'h6)] ^~ $unsigned(reg525))} : reg559) ?
                  reg452 : {(wire449[(4'ha):(4'ha)] * reg546)});
              reg575 = reg559[(1'h0):(1'h0)];
            end
          else
            begin
              reg576 <= $unsigned((~&$unsigned((-reg572))));
              reg577 = forvar572;
            end
          reg578 = $signed(reg457[(4'hc):(3'h6)]);
          for (forvar579 = (1'h0); (forvar579 < (1'h1)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 = $signed(reg541);
              reg581 = (({$signed(reg472)} > $signed($signed(((8'ha6) >= reg552)))) > ((($signed(reg459) == (reg518 ?
                          reg473 : reg568)) ?
                      $unsigned($signed((8'hb5))) : reg580) ?
                  reg461 : $unsigned($signed(((8'hbb) | reg571)))));
              reg582 <= reg536[(2'h3):(2'h3)];
              reg583 <= (~&{{$signed($unsigned(reg531))},
                  (((reg488 >>> reg510) ?
                          (!reg549) : (reg500 ? reg494 : reg525)) ?
                      $signed(reg464) : reg527[(1'h1):(1'h1)])});
            end
          if (wire563[(2'h3):(1'h1)])
            begin
              reg584 = ((($signed(reg503) && ($unsigned((8'hba)) ?
                      reg583 : (reg567 ^~ reg566))) ?
                  reg452[(3'h6):(3'h4)] : (-reg567[(4'hf):(4'hb)])) == reg502);
            end
          else
            begin
              reg584 = reg466;
              reg585 = $unsigned(forvar579[(3'h6):(2'h3)]);
              reg586 <= ({wire449,
                      $signed($unsigned((reg503 ? wire564 : reg494)))} ?
                  reg550 : {reg572});
            end
        end
    end
  assign wire587 = $unsigned($unsigned($unsigned((^~reg582[(3'h6):(3'h5)]))));
  always
    @(posedge clk) begin
      if ($signed({$unsigned(($unsigned(reg536) & (reg549 ?
              reg486 : reg559)))}))
        begin
          for (forvar588 = (1'h0); (forvar588 < (1'h1)); forvar588 = (forvar588 + (1'h1)))
            begin
              reg589 = (~|$signed($unsigned((!(|(8'ha0))))));
              reg590 <= (8'hb0);
              reg591 <= wire450[(4'he):(1'h1)];
            end
          if ($unsigned($signed(wire561)))
            begin
              reg592 <= (~&reg505);
              reg593 = {{($signed(reg558) << (|wire564))}};
              reg594 <= ((!reg590[(3'h6):(3'h4)]) > $unsigned($signed((+reg479[(4'hc):(4'hc)]))));
              reg595 = reg466[(2'h2):(2'h2)];
            end
          else
            begin
              reg593 = $signed((~reg524[(2'h3):(2'h3)]));
            end
          for (forvar596 = (1'h0); (forvar596 < (3'h4)); forvar596 = (forvar596 + (1'h1)))
            begin
              reg597 <= $signed(((wire450[(5'h10):(4'hd)] && $signed((reg506 ?
                      reg547 : reg488))) ?
                  (8'hb2) : reg510[(1'h0):(1'h0)]));
              reg598 = ($signed(($unsigned((wire561 ? reg569 : forvar596)) ?
                      (reg538 ?
                          (8'hb5) : $signed((8'h9e))) : $unsigned((~^reg466)))) ?
                  ($unsigned($signed(((8'hae) ?
                      reg472 : reg582))) >> (reg486[(4'h9):(2'h3)] ?
                      $unsigned($unsigned((8'h9c))) : (^(reg567 ?
                          (8'h9c) : reg472)))) : (^(-(reg552 - wire450[(3'h4):(1'h0)]))));
            end
          reg599 = {$unsigned($signed($unsigned(reg583)))};
        end
      else
        begin
          reg588 <= reg467;
          reg590 <= reg542[(4'hd):(4'hb)];
          reg591 <= $unsigned($signed(reg538));
          reg592 <= reg542[(4'h8):(3'h7)];
          reg594 <= reg483[(2'h2):(2'h2)];
        end
      if ((+$unsigned(((wire561 * (|reg538)) ?
          (reg576[(4'hb):(3'h6)] + (wire562 ~^ reg520)) : wire563[(3'h5):(2'h2)]))))
        begin
          if (((wire562 ?
              {$signed($unsigned(reg500))} : $signed(reg524[(3'h6):(2'h3)])) <= $signed(reg500)))
            begin
              reg600 = (!$unsigned(reg583[(3'h6):(3'h5)]));
              reg601 <= ((~&$signed($unsigned($unsigned((8'hb6))))) ?
                  $unsigned({$unsigned((reg572 << reg466)),
                      $signed(reg506)}) : reg457[(2'h3):(2'h3)]);
            end
          else
            begin
              reg600 = $signed(reg526);
            end
          if (reg486)
            begin
              reg602 = ((~^$unsigned(reg466)) ~^ ($signed((+(wire448 | reg483))) - reg461));
              reg603 <= (~&(reg525[(4'hf):(4'ha)] ?
                  $signed(reg510[(3'h6):(2'h2)]) : ($unsigned(reg598[(4'hb):(3'h4)]) ?
                      (~|{reg597, wire561}) : (!$unsigned(reg556)))));
              reg604 <= (reg590[(3'h4):(1'h1)] <<< reg488);
              reg605 = (reg567[(5'h15):(4'hd)] - $signed((~^(reg486 ?
                  (reg472 ? reg603 : reg589) : $signed(reg464)))));
              reg606 <= reg503[(2'h2):(2'h2)];
            end
          else
            begin
              reg602 = $unsigned({($unsigned($signed(reg546)) < wire564)});
              reg605 = {(reg576 - reg549[(1'h1):(1'h0)])};
            end
        end
      else
        begin
          if ($signed(((^(~$signed(wire449))) <<< (reg600[(2'h2):(1'h1)] ?
              (reg565[(2'h2):(1'h1)] ?
                  (!reg598) : (wire561 < reg602)) : $unsigned(((8'hb5) + reg525))))))
            begin
              reg601 <= reg466;
              reg602 = reg473[(4'hb):(3'h7)];
              reg603 <= ({(^((reg480 <= reg571) || (reg488 ?
                          reg565 : reg558)))} ?
                  {reg590} : ({reg489[(2'h2):(2'h2)]} | $unsigned(reg602)));
            end
          else
            begin
              reg601 <= reg506[(3'h4):(1'h0)];
              reg603 <= ({$unsigned((^~$unsigned(reg552))),
                  (reg604 ?
                      wire450[(4'hb):(2'h3)] : $signed(reg550))} <= (reg525[(4'hf):(4'h9)] >>> (reg538[(3'h4):(3'h4)] ?
                  $unsigned(reg520) : (|$signed(reg591)))));
            end
          for (forvar604 = (1'h0); (forvar604 < (2'h3)); forvar604 = (forvar604 + (1'h1)))
            begin
              reg605 = ($unsigned(($unsigned((reg589 >> reg532)) <= reg503[(2'h3):(1'h0)])) >>> reg598);
              reg606 <= {(8'hb9), (~&(^~wire561))};
              reg607 <= $unsigned(wire564[(1'h1):(1'h0)]);
            end
          for (forvar608 = (1'h0); (forvar608 < (1'h0)); forvar608 = (forvar608 + (1'h1)))
            begin
              reg609 <= $signed($signed(reg455[(1'h1):(1'h1)]));
              reg610 <= reg583;
              reg611 <= ($unsigned((($unsigned(reg601) ?
                          (reg532 ?
                              reg583 : reg571) : reg609[(5'h14):(5'h13)]) ?
                      ($unsigned(wire587) <<< reg531[(1'h1):(1'h0)]) : {(^wire563)})) ?
                  (reg605[(1'h1):(1'h0)] ?
                      (8'had) : (reg527[(4'hf):(4'h8)] ?
                          ((~reg486) ?
                              (reg513 ? reg605 : reg510) : {reg586,
                                  (7'h42)}) : {reg547})) : reg489);
              reg612 <= reg520[(4'he):(3'h4)];
              reg613 <= ((8'hbe) ?
                  (~&(($unsigned(reg588) ?
                          ((8'ha2) ? reg595 : wire561) : $unsigned(reg457)) ?
                      reg492 : (^~$unsigned(reg549)))) : $signed($unsigned({$signed(wire450)})));
            end
        end
      reg614 = reg590;
      reg615 <= (reg592 >> (8'ha9));
    end
  assign wire616 = $signed(reg603[(1'h1):(1'h0)]);
  assign wire617 = $unsigned(reg550[(3'h5):(1'h1)]);
  assign wire618 = (&$signed((~&({reg552} >> (wire447 ? wire563 : reg467)))));
  always
    @(posedge clk) begin
      if ((8'hbf))
        begin
          if ((!$unsigned($signed($signed(reg455[(3'h5):(2'h3)])))))
            begin
              reg619 <= (!(reg594[(4'h8):(1'h0)] && $signed((reg488 & (~|(8'ha1))))));
              reg620 <= $signed(reg467);
              reg621 = reg489[(1'h1):(1'h0)];
            end
          else
            begin
              reg621 = ($signed(reg615[(4'hc):(4'h8)]) ?
                  ($unsigned(($unsigned(wire561) > reg591[(4'ha):(3'h7)])) ?
                      reg455[(1'h0):(1'h0)] : $unsigned((|(reg559 ?
                          reg526 : reg503)))) : reg527[(5'h15):(3'h5)]);
              reg622 = $unsigned((^~{reg500[(3'h4):(1'h1)]}));
              reg623 <= $signed(reg615);
              reg624 <= $unsigned(reg594[(4'h9):(2'h2)]);
              reg625 <= $unsigned($signed(((^reg601) ?
                  reg610 : {(reg588 & (8'h9e)), (reg532 ? wire447 : reg489)})));
            end
          reg626 = (^~{reg536[(3'h4):(3'h4)]});
          for (forvar627 = (1'h0); (forvar627 < (2'h3)); forvar627 = (forvar627 + (1'h1)))
            begin
              reg628 = ((($unsigned($unsigned(wire564)) ?
                      reg502 : ($signed(wire564) + $signed(reg569))) <= wire447) ?
                  (forvar627 ?
                      ((wire560 ? reg538[(4'h8):(2'h3)] : $signed(reg518)) ?
                          $signed((wire560 ?
                              reg518 : forvar627)) : $unsigned($unsigned(wire447))) : (!(7'h46))) : reg606[(2'h2):(1'h0)]);
              reg629 = ((reg559 ?
                  reg601[(1'h0):(1'h0)] : $signed({(8'had)})) & reg526);
              reg630 <= ($signed((-reg518)) && reg571[(5'h11):(4'hf)]);
              reg631 <= $signed(wire449);
              reg632 = reg527[(3'h5):(1'h0)];
            end
        end
      else
        begin
          reg621 = $unsigned(($unsigned($unsigned((forvar627 | reg527))) ?
              reg613 : reg456[(2'h3):(1'h0)]));
        end
      for (forvar633 = (1'h0); (forvar633 < (2'h2)); forvar633 = (forvar633 + (1'h1)))
        begin
          reg634 <= $unsigned(($signed({(~reg613)}) >= (^~((reg590 ?
                  reg572 : forvar633) ?
              (!reg455) : reg597))));
          for (forvar635 = (1'h0); (forvar635 < (1'h0)); forvar635 = (forvar635 + (1'h1)))
            begin
              reg636 = (reg557[(2'h2):(2'h2)] ?
                  (~($signed((wire617 | reg604)) ?
                      $signed($signed(reg477)) : {$unsigned(reg467)})) : (+($unsigned((reg626 ?
                          wire448 : reg536)) ?
                      reg526[(3'h5):(3'h5)] : ((reg473 >= reg466) <= $signed((8'hb6))))));
            end
          reg637 <= $unsigned($unsigned($unsigned(reg455[(2'h2):(1'h1)])));
          if (reg456[(1'h0):(1'h0)])
            begin
              reg638 <= {(reg603 ?
                      (~$unsigned((reg538 & (7'h46)))) : reg538[(3'h5):(2'h2)]),
                  reg503[(3'h4):(1'h1)]};
            end
          else
            begin
              reg638 <= (^({$signed(reg467[(2'h2):(1'h0)]),
                  ((wire618 <= reg524) ? reg606 : reg565)} - {{(^reg612)}}));
              reg639 <= (^~($signed(($unsigned(reg610) ?
                      $unsigned(reg538) : $unsigned((8'hbe)))) ?
                  (reg547 ?
                      ((wire450 ?
                          reg500 : reg591) <<< $signed((8'had))) : $signed($signed(wire617))) : $signed($signed($unsigned(reg567)))));
              reg640 = (reg591[(1'h1):(1'h0)] >= (-$signed((reg571 >= reg565[(1'h1):(1'h1)]))));
              reg641 <= reg557;
              reg642 = $signed((reg620[(4'hb):(4'h9)] + reg488));
            end
        end
    end
  assign wire643 = (8'hab);
  always
    @(posedge clk) begin
      reg644 <= ($signed((reg611[(2'h3):(2'h3)] == $unsigned({reg547,
              wire617}))) ?
          wire449[(4'hc):(3'h6)] : reg586[(3'h5):(2'h3)]);
    end
  assign wire645 = $signed(reg503[(2'h3):(1'h0)]);
  assign wire646 = $unsigned({$signed(($signed(reg556) ?
                           (|reg597) : (reg603 << wire587)))});
  always
    @(posedge clk) begin
      if (wire645[(2'h2):(1'h1)])
        begin
          reg647 = ({$unsigned({$signed((8'haf))}),
                  {({reg549, reg542} & $unsigned(reg486)),
                      $unsigned({reg504})}} ?
              ((((8'hb0) >>> (~(8'hae))) * (reg572[(3'h7):(3'h6)] | $unsigned(reg546))) ?
                  (((reg531 ? reg472 : reg606) ?
                      $signed(reg452) : $signed(reg637)) >= reg559) : (((!wire587) ?
                      {reg644} : (-reg541)) != {(~^reg483)})) : wire618);
          reg648 <= reg524;
        end
      else
        begin
          reg648 <= $unsigned((~(((reg601 != reg477) <<< (wire561 == wire645)) ?
              reg594[(4'h8):(3'h4)] : ($unsigned(wire560) > reg606))));
          for (forvar649 = (1'h0); (forvar649 < (2'h3)); forvar649 = (forvar649 + (1'h1)))
            begin
              reg650 = reg457;
              reg651 <= (((reg526 ? reg604[(3'h4):(3'h4)] : reg592) ?
                      $signed(reg473[(4'hd):(2'h2)]) : ($unsigned(((8'ha9) ?
                              reg505 : (8'hb7))) ?
                          $signed(reg526) : $unsigned((reg588 == reg625)))) ?
                  $signed((+(7'h44))) : ($signed($signed(reg630)) ?
                      reg606 : reg623));
            end
          for (forvar652 = (1'h0); (forvar652 < (2'h2)); forvar652 = (forvar652 + (1'h1)))
            begin
              reg653 <= (($unsigned(($unsigned(reg525) && wire646[(3'h5):(2'h3)])) > $unsigned((~&(reg538 && reg611)))) ^~ reg647);
              reg654 = {($unsigned(((8'h9c) ?
                          (&reg624) : (wire645 ? reg541 : reg502))) ?
                      (((^~reg492) + $signed(forvar649)) ?
                          reg513 : ((^~reg456) ?
                              reg527 : (reg647 == reg653))) : (((reg620 ?
                                  reg494 : reg606) ?
                              (reg455 ? (7'h45) : wire561) : ((7'h41) ?
                                  reg582 : wire449)) ?
                          (^~reg543[(4'hb):(4'hb)]) : reg588)),
                  $unsigned(wire587[(3'h4):(2'h2)])};
              reg655 = ((+(($unsigned(reg473) <= $signed(reg631)) ?
                      (reg459[(2'h2):(1'h0)] || (reg592 <<< reg531)) : $signed((wire618 != reg653)))) ?
                  (!($signed((wire617 ? wire561 : reg488)) ?
                      ((reg610 ? reg631 : (7'h41)) ?
                          reg525 : (reg653 ?
                              reg576 : reg455)) : reg588[(4'hf):(4'h9)])) : $unsigned(($unsigned(((7'h46) ?
                          reg569 : reg620)) ?
                      (^(reg567 | (8'hbe))) : (~^reg507))));
              reg656 = (8'ha7);
            end
          reg657 <= $unsigned((reg615[(1'h0):(1'h0)] ?
              $unsigned(reg582) : forvar649[(1'h1):(1'h0)]));
        end
    end
  assign wire658 = $signed((!({(reg541 ^ reg483)} ?
                       (~&reg648[(5'h12):(2'h2)]) : reg546[(3'h4):(1'h0)])));
  assign wire659 = {reg542};
  always
    @(posedge clk) begin
      reg660 = {reg531, $signed((reg639 >>> (~(reg624 - reg524))))};
      for (forvar661 = (1'h0); (forvar661 < (2'h2)); forvar661 = (forvar661 + (1'h1)))
        begin
          for (forvar662 = (1'h0); (forvar662 < (2'h3)); forvar662 = (forvar662 + (1'h1)))
            begin
              reg663 = $signed(((~reg532) > reg653));
              reg664 = reg479[(2'h3):(1'h1)];
              reg665 <= (8'hab);
            end
        end
      reg666 <= ($signed($signed(reg639)) ?
          (reg572[(1'h0):(1'h0)] ?
              reg592 : (|$signed($signed(reg518)))) : (-(8'hb8)));
      reg667 <= ($unsigned(reg606[(4'h8):(3'h6)]) ^~ {(~^{(-(7'h43))})});
      for (forvar668 = (1'h0); (forvar668 < (1'h0)); forvar668 = (forvar668 + (1'h1)))
        begin
          reg669 = $signed(({wire617} >>> ({reg506} & (^$unsigned(reg461)))));
          reg670 <= ($unsigned((reg603 ?
                  reg550[(3'h6):(3'h5)] : (|$unsigned(reg538)))) ?
              (-reg507[(3'h5):(3'h5)]) : $signed((^~(7'h40))));
          for (forvar671 = (1'h0); (forvar671 < (3'h4)); forvar671 = (forvar671 + (1'h1)))
            begin
              reg672 = $signed(wire564);
              reg673 <= reg541[(2'h2):(1'h1)];
            end
          reg674 <= ($signed((8'ha8)) >> $signed((-(wire616[(3'h6):(3'h4)] <<< (reg612 >>> reg613)))));
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed((~|$unsigned({reg531, reg486})))))
        begin
          if ((~$signed(reg639[(1'h0):(1'h0)])))
            begin
              reg675 = $unsigned($unsigned($signed((reg531[(1'h1):(1'h0)] != $unsigned(reg591)))));
              reg676 = wire616[(3'h4):(2'h2)];
              reg677 = reg525;
              reg678 <= (8'ha4);
              reg679 = reg597;
            end
          else
            begin
              reg675 = $signed(wire564[(3'h4):(2'h3)]);
              reg678 <= ($unsigned($unsigned(reg648[(4'h8):(2'h3)])) != {wire564[(4'hb):(2'h3)],
                  $signed(reg503)});
              reg680 <= $unsigned((reg571[(5'h12):(4'he)] ?
                  reg507[(4'h9):(3'h5)] : ($unsigned((reg653 | reg525)) ?
                      {((8'hbe) ? reg461 : reg455),
                          (~reg510)} : (-$unsigned(reg520)))));
            end
          for (forvar681 = (1'h0); (forvar681 < (3'h4)); forvar681 = (forvar681 + (1'h1)))
            begin
              reg682 = $signed($signed(((-$signed(reg565)) >= $signed((wire618 ?
                  reg503 : (7'h43))))));
            end
          for (forvar683 = (1'h0); (forvar683 < (2'h3)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 <= (reg504[(4'hc):(1'h1)] ^~ {((reg549 << (^reg489)) != {reg601[(2'h3):(2'h3)]}),
                  ($signed({reg556, reg641}) ?
                      (~|reg607[(2'h3):(2'h2)]) : reg682)});
              reg685 <= $unsigned(($unsigned($unsigned((~&reg557))) << ({reg576,
                  (8'h9d)} ~^ $signed(reg494[(3'h7):(1'h0)]))));
            end
          if ({(8'h9c)})
            begin
              reg686 = $unsigned((^($signed((~^(8'hb3))) ?
                  reg680[(5'h15):(5'h14)] : (((8'hb3) ? wire646 : (8'hb0)) ?
                      (-reg506) : reg486))));
              reg687 = $signed(reg679[(3'h7):(3'h6)]);
              reg688 <= (+{reg558[(5'h16):(3'h6)]});
              reg689 = $unsigned(reg506);
            end
          else
            begin
              reg688 <= (reg688[(2'h2):(2'h2)] <= reg524[(3'h5):(3'h4)]);
              reg689 = ((^~reg473) << $unsigned((reg510 ?
                  ((reg677 ? reg510 : reg592) ~^ reg592) : reg536)));
              reg690 <= reg467;
              reg691 <= ($signed(reg619) ?
                  reg464[(4'ha):(3'h5)] : ($signed(reg666[(4'he):(2'h3)]) ?
                      ((^(reg538 ~^ reg637)) ?
                          ((reg657 >>> (8'hab)) ?
                              $unsigned(reg510) : (reg674 ?
                                  reg452 : reg673)) : reg459) : (((reg685 ?
                              reg505 : reg565) ?
                          reg480 : $signed(reg610)) ^ (wire448 ?
                          wire587[(3'h5):(3'h5)] : reg571[(5'h11):(4'ha)]))));
            end
          for (forvar692 = (1'h0); (forvar692 < (2'h3)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 <= ((8'hb6) <= (8'h9f));
            end
        end
      else
        begin
          for (forvar675 = (1'h0); (forvar675 < (1'h1)); forvar675 = (forvar675 + (1'h1)))
            begin
              reg678 <= $signed({reg572[(3'h7):(3'h4)],
                  ($signed($signed(wire587)) ?
                      reg518[(1'h1):(1'h0)] : (~|$unsigned((8'ha2))))});
            end
          for (forvar679 = (1'h0); (forvar679 < (1'h0)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 <= $unsigned($unsigned(reg687));
              reg681 <= reg467[(5'h10):(4'h9)];
              reg682 = (($unsigned({$unsigned(reg624)}) <<< {{(reg677 ?
                          reg673 : reg634)},
                  {(^~reg504),
                      reg631}}) == $signed($unsigned(reg680[(4'hb):(3'h4)])));
              reg683 <= {(&forvar681[(4'h9):(4'h9)])};
              reg686 = $unsigned({reg459, (^wire563)});
            end
          reg688 <= {reg615[(1'h1):(1'h0)], reg507[(3'h4):(2'h2)]};
          reg690 <= ($signed((~({reg675, reg510} ?
              reg510[(2'h2):(2'h2)] : reg556[(4'hf):(4'h8)]))) >>> (((((8'hab) != reg683) ?
              {reg603, reg588} : {reg693,
                  (8'hae)}) > $unsigned(wire561)) && (&{reg556[(2'h3):(1'h0)],
              (reg588 ? reg559 : reg583)})));
          if ($signed(wire560))
            begin
              reg692 = reg592;
              reg693 <= (~$unsigned((reg456[(1'h1):(1'h1)] ?
                  ($unsigned(wire447) ?
                      $unsigned(reg639) : $signed((8'ha2))) : $signed(reg644))));
            end
          else
            begin
              reg692 = reg597[(2'h2):(2'h2)];
            end
        end
    end
endmodule
(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'haa5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire0;
  input wire [(5'h12):(1'h0)] wire1;
  input wire signed [(4'hd):(1'h0)] wire2;
  input wire [(5'h14):(1'h0)] wire3;
  input wire [(4'h9):(1'h0)] wire4;
  reg [(5'h13):(1'h0)] reg958 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg957 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg956 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar955 = (1'h0);
  reg [(4'h8):(1'h0)] reg954 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg953 = (1'h0);
  reg [(5'h13):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg951 = (1'h0);
  reg [(5'h15):(1'h0)] reg950 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg948 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg946 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg945 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar944 = (1'h0);
  reg [(3'h6):(1'h0)] forvar943 = (1'h0);
  reg [(2'h3):(1'h0)] reg942 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg941 = (1'h0);
  reg [(5'h13):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg939 = (1'h0);
  reg [(4'hd):(1'h0)] reg938 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar937 = (1'h0);
  reg [(4'hf):(1'h0)] reg925 = (1'h0);
  reg [(5'h14):(1'h0)] forvar923 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg936 = (1'h0);
  reg [(2'h3):(1'h0)] reg935 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar934 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg933 = (1'h0);
  reg [(3'h4):(1'h0)] reg932 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg931 = (1'h0);
  reg [(4'h8):(1'h0)] forvar930 = (1'h0);
  reg [(5'h15):(1'h0)] reg929 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg928 = (1'h0);
  reg [(5'h15):(1'h0)] reg927 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg926 = (1'h0);
  reg [(4'hf):(1'h0)] forvar925 = (1'h0);
  reg [(4'hf):(1'h0)] reg924 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg923 = (1'h0);
  reg [(4'hd):(1'h0)] reg922 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg921 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg920 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar919 = (1'h0);
  reg [(2'h3):(1'h0)] reg918 = (1'h0);
  reg [(5'h10):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg916 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg915 = (1'h0);
  reg [(5'h11):(1'h0)] forvar914 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire882;
  reg [(5'h11):(1'h0)] reg881 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar879 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg878 = (1'h0);
  reg [(5'h15):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg876 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg875 = (1'h0);
  reg [(4'he):(1'h0)] forvar874 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg873 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg872 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg871 = (1'h0);
  reg [(5'h14):(1'h0)] reg870 = (1'h0);
  reg [(4'ha):(1'h0)] forvar869 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg868 = (1'h0);
  reg [(5'h11):(1'h0)] forvar867 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar866 = (1'h0);
  reg [(3'h5):(1'h0)] reg865 = (1'h0);
  reg [(5'h12):(1'h0)] reg864 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg863 = (1'h0);
  reg [(3'h7):(1'h0)] reg862 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg861 = (1'h0);
  reg [(3'h5):(1'h0)] forvar860 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg859 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar858 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg852 = (1'h0);
  reg [(5'h10):(1'h0)] forvar851 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg846 = (1'h0);
  reg [(3'h6):(1'h0)] forvar845 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg857 = (1'h0);
  reg signed [(4'he):(1'h0)] reg856 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg854 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg853 = (1'h0);
  reg [(5'h12):(1'h0)] forvar852 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg850 = (1'h0);
  reg [(4'hd):(1'h0)] reg849 = (1'h0);
  reg [(4'h9):(1'h0)] reg848 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar846 = (1'h0);
  reg [(3'h5):(1'h0)] reg845 = (1'h0);
  reg [(2'h3):(1'h0)] reg844 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire5;
  wire signed [(4'hd):(1'h0)] wire6;
  wire signed [(5'h13):(1'h0)] wire7;
  reg signed [(5'h11):(1'h0)] forvar8 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg9 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar10 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg12 = (1'h0);
  reg [(4'h9):(1'h0)] forvar13 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar14 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg15 = (1'h0);
  reg [(4'ha):(1'h0)] reg16 = (1'h0);
  reg [(5'h13):(1'h0)] reg17 = (1'h0);
  reg [(4'hb):(1'h0)] forvar18 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar19 = (1'h0);
  reg [(5'h15):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg21 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg22 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar23 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg24 = (1'h0);
  reg [(5'h11):(1'h0)] reg25 = (1'h0);
  reg [(4'he):(1'h0)] forvar26 = (1'h0);
  reg [(5'h11):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg28 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg29 = (1'h0);
  reg [(2'h3):(1'h0)] reg30 = (1'h0);
  reg [(2'h2):(1'h0)] reg31 = (1'h0);
  reg [(5'h11):(1'h0)] reg32 = (1'h0);
  reg [(5'h10):(1'h0)] reg33 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg34 = (1'h0);
  reg [(4'hf):(1'h0)] reg35 = (1'h0);
  reg [(5'h10):(1'h0)] reg36 = (1'h0);
  reg [(2'h3):(1'h0)] reg37 = (1'h0);
  reg [(3'h7):(1'h0)] forvar38 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar39 = (1'h0);
  reg [(3'h5):(1'h0)] reg40 = (1'h0);
  reg [(4'he):(1'h0)] reg41 = (1'h0);
  reg [(5'h15):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg43 = (1'h0);
  reg [(5'h11):(1'h0)] reg44 = (1'h0);
  reg [(5'h10):(1'h0)] forvar45 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg48 = (1'h0);
  reg [(2'h3):(1'h0)] reg49 = (1'h0);
  reg [(2'h2):(1'h0)] reg50 = (1'h0);
  wire [(4'he):(1'h0)] wire557;
  wire signed [(5'h14):(1'h0)] wire559;
  wire [(5'h10):(1'h0)] wire560;
  wire [(4'h9):(1'h0)] wire561;
  reg [(4'hb):(1'h0)] reg562 = (1'h0);
  reg [(4'hd):(1'h0)] reg563 = (1'h0);
  reg [(4'hd):(1'h0)] reg564 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar562 = (1'h0);
  reg [(4'hd):(1'h0)] forvar565 = (1'h0);
  reg [(3'h7):(1'h0)] reg566 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar567 = (1'h0);
  reg [(5'h15):(1'h0)] reg568 = (1'h0);
  reg [(3'h4):(1'h0)] reg569 = (1'h0);
  reg [(4'hd):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar572 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg573 = (1'h0);
  reg [(4'hc):(1'h0)] reg574 = (1'h0);
  reg [(4'hf):(1'h0)] reg575 = (1'h0);
  reg [(5'h15):(1'h0)] reg576 = (1'h0);
  reg [(4'hc):(1'h0)] reg577 = (1'h0);
  reg [(4'ha):(1'h0)] forvar578 = (1'h0);
  reg [(4'h9):(1'h0)] reg579 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg581 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg582 = (1'h0);
  reg [(5'h10):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg584 = (1'h0);
  reg [(4'hf):(1'h0)] reg578 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar582 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg585 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg586 = (1'h0);
  reg [(4'hc):(1'h0)] reg587 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar588 = (1'h0);
  reg [(5'h13):(1'h0)] reg589 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar592 = (1'h0);
  reg signed [(4'he):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar595 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg596 = (1'h0);
  reg [(5'h11):(1'h0)] reg597 = (1'h0);
  reg [(2'h3):(1'h0)] reg598 = (1'h0);
  reg [(5'h10):(1'h0)] reg599 = (1'h0);
  reg [(4'h9):(1'h0)] reg600 = (1'h0);
  reg [(3'h5):(1'h0)] reg601 = (1'h0);
  reg [(3'h7):(1'h0)] forvar602 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar603 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg605 = (1'h0);
  reg [(3'h6):(1'h0)] reg606 = (1'h0);
  reg [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar608 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg609 = (1'h0);
  reg [(5'h10):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar611 = (1'h0);
  reg [(4'he):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg613 = (1'h0);
  reg [(4'hb):(1'h0)] reg614 = (1'h0);
  wire [(4'hf):(1'h0)] wire842;
  reg [(3'h5):(1'h0)] forvar884 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg885 = (1'h0);
  reg [(4'h8):(1'h0)] forvar886 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg887 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg888 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg889 = (1'h0);
  reg [(5'h10):(1'h0)] reg890 = (1'h0);
  reg [(5'h15):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar892 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg893 = (1'h0);
  reg [(3'h6):(1'h0)] reg894 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg895 = (1'h0);
  reg [(5'h12):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg897 = (1'h0);
  reg [(4'hf):(1'h0)] reg898 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar899 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar900 = (1'h0);
  reg [(5'h13):(1'h0)] reg901 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg902 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg903 = (1'h0);
  reg [(5'h11):(1'h0)] forvar904 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg905 = (1'h0);
  reg [(5'h14):(1'h0)] reg906 = (1'h0);
  reg [(4'he):(1'h0)] reg907 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire908;
  wire signed [(4'hb):(1'h0)] wire909;
  wire signed [(2'h2):(1'h0)] wire910;
  wire [(5'h14):(1'h0)] wire911;
  wire [(5'h12):(1'h0)] wire912;
  assign y = {reg958,
                 reg957,
                 reg956,
                 forvar955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 reg945,
                 forvar944,
                 forvar943,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg925,
                 forvar923,
                 reg919,
                 reg936,
                 reg935,
                 forvar934,
                 reg933,
                 reg932,
                 reg931,
                 forvar930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 forvar925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 forvar919,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 forvar914,
                 wire882,
                 reg881,
                 reg880,
                 forvar879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 forvar874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 forvar869,
                 reg868,
                 forvar867,
                 forvar866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 forvar860,
                 reg859,
                 forvar858,
                 reg852,
                 forvar851,
                 reg846,
                 forvar845,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 forvar852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 forvar846,
                 reg845,
                 reg844,
                 wire5,
                 wire6,
                 wire7,
                 forvar8,
                 reg9,
                 forvar10,
                 reg11,
                 reg12,
                 forvar13,
                 forvar14,
                 reg15,
                 reg16,
                 reg17,
                 forvar18,
                 forvar19,
                 reg20,
                 reg21,
                 reg22,
                 forvar23,
                 reg24,
                 reg25,
                 forvar26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 forvar38,
                 forvar39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 forvar45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 wire557,
                 wire559,
                 wire560,
                 wire561,
                 reg562,
                 reg563,
                 reg564,
                 forvar562,
                 forvar565,
                 reg566,
                 forvar567,
                 reg568,
                 reg569,
                 reg570,
                 reg571,
                 forvar572,
                 reg573,
                 reg574,
                 reg575,
                 reg576,
                 reg577,
                 forvar578,
                 reg579,
                 reg580,
                 reg581,
                 reg582,
                 reg583,
                 reg584,
                 reg578,
                 forvar582,
                 reg585,
                 reg586,
                 reg587,
                 forvar588,
                 reg589,
                 reg590,
                 reg591,
                 forvar592,
                 reg593,
                 reg594,
                 forvar595,
                 reg596,
                 reg597,
                 reg598,
                 reg599,
                 reg600,
                 reg601,
                 forvar602,
                 forvar603,
                 reg604,
                 reg605,
                 reg606,
                 reg607,
                 forvar608,
                 reg609,
                 reg610,
                 forvar611,
                 reg612,
                 reg613,
                 reg614,
                 wire842,
                 forvar884,
                 reg885,
                 forvar886,
                 reg887,
                 reg888,
                 reg889,
                 reg890,
                 reg891,
                 forvar892,
                 reg893,
                 reg894,
                 reg895,
                 reg896,
                 reg897,
                 reg898,
                 forvar899,
                 forvar900,
                 reg901,
                 reg902,
                 reg903,
                 forvar904,
                 reg905,
                 reg906,
                 reg907,
                 wire908,
                 wire909,
                 wire910,
                 wire911,
                 wire912,
                 (1'h0)};
  assign wire5 = $unsigned($signed($signed(($signed(wire1) <<< $unsigned((7'h41))))));
  assign wire6 = (-wire2[(3'h7):(2'h2)]);
  assign wire7 = {$signed(wire4),
                     (((~wire2) >> wire4) && $signed((~^wire2[(3'h7):(1'h1)])))};
  always
    @(posedge clk) begin
      for (forvar8 = (1'h0); (forvar8 < (1'h1)); forvar8 = (forvar8 + (1'h1)))
        begin
          reg9 <= (((8'hac) ? (7'h41) : $signed(wire2)) ?
              (wire4 ^ (~|$unsigned($signed(forvar8)))) : $signed(((8'ha6) | wire5[(2'h2):(1'h1)])));
          for (forvar10 = (1'h0); (forvar10 < (2'h2)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 = wire5;
              reg12 = {{$unsigned(forvar10[(1'h1):(1'h1)])},
                  {wire0[(4'h8):(1'h0)],
                      (wire2[(4'hb):(3'h4)] ?
                          $signed(((8'hbd) | reg9)) : $unsigned($signed((8'h9e))))}};
            end
        end
      for (forvar13 = (1'h0); (forvar13 < (2'h3)); forvar13 = (forvar13 + (1'h1)))
        begin
          for (forvar14 = (1'h0); (forvar14 < (1'h0)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= (wire2 * (|{{$signed(forvar10), wire5[(3'h5):(1'h1)]}}));
            end
          reg16 <= {reg11[(1'h1):(1'h0)]};
        end
      reg17 = reg9;
    end
  always
    @(posedge clk) begin
      for (forvar18 = (1'h0); (forvar18 < (1'h0)); forvar18 = (forvar18 + (1'h1)))
        begin
          for (forvar19 = (1'h0); (forvar19 < (2'h3)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 <= wire5;
              reg21 <= $signed("hcmb3gMxq4");
              reg22 <= "qyVrc9QBTKwH";
            end
          for (forvar23 = (1'h0); (forvar23 < (3'h4)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 <= ((-{((wire7 ? forvar8 : reg15) ?
                      $signed(wire7) : (reg9 <<< reg17)),
                  ({reg15,
                      (8'h9d)} <<< (8'ha1))}) != (~^{($unsigned(forvar14) != (8'hbd))}));
              reg25 <= reg24;
            end
          for (forvar26 = (1'h0); (forvar26 < (2'h3)); forvar26 = (forvar26 + (1'h1)))
            begin
              reg27 <= (8'ha8);
              reg28 <= ($signed(wire2) ?
                  $unsigned((((~&forvar19) | $signed(forvar18)) ?
                      reg25[(4'he):(4'hd)] : (&$signed(wire1)))) : (^~(^~(^{(8'hae),
                      wire0}))));
            end
          if ($unsigned(reg17[(1'h1):(1'h1)]))
            begin
              reg29 <= {wire3[(5'h11):(3'h6)]};
              reg30 = reg29;
              reg31 = ($unsigned(wire5) != reg20);
              reg32 <= $signed($signed((^~{((8'hbd) << reg12)})));
              reg33 <= ((~|(forvar19[(3'h4):(1'h1)] > (reg22[(2'h2):(1'h0)] ?
                      (-forvar19) : ((8'hb3) & forvar18)))) ?
                  $unsigned(forvar26) : $signed(((-(reg25 ^ reg11)) ?
                      $unsigned(((8'hb1) ? wire3 : (8'ha8))) : reg22)));
            end
          else
            begin
              reg29 = reg20;
              reg30 <= (({{(reg12 ? reg33 : forvar14), $unsigned(reg31)}} ?
                  $unsigned(reg31) : (^~({(8'hb3), reg28} ?
                      "pb0DDU320sLpAoz3LLR" : (reg22 ?
                          reg16 : wire3)))) & forvar13);
              reg31 <= (-(8'hbc));
              reg32 = {$unsigned(reg11),
                  (~^$signed(((wire4 ? reg12 : reg29) ~^ (forvar23 > reg21))))};
            end
          if (reg33)
            begin
              reg34 = {($unsigned(reg9[(3'h7):(2'h2)]) ?
                      (~^$signed("wwCrZx8C")) : {(reg21 ?
                              (reg24 ? reg15 : wire7) : wire0[(1'h1):(1'h1)])}),
                  ("mzWBr2QYAuLt" ?
                      (~$signed(wire2[(1'h0):(1'h0)])) : (~^$signed($signed((8'h9d)))))};
              reg35 <= (&reg33);
              reg36 = {(reg24 == {(~&reg31[(1'h0):(1'h0)])}), forvar26};
              reg37 = ($signed(forvar13[(1'h0):(1'h0)]) ?
                  $signed(reg25) : $signed($unsigned(($signed((7'h43)) ?
                      (+forvar23) : (!reg21)))));
            end
          else
            begin
              reg34 = forvar8;
              reg35 = ((^~forvar19[(1'h0):(1'h0)]) ?
                  (-(forvar8 ?
                      {(8'hbc),
                          reg9} : "9Wi1YSxwSpGEi")) : (((-(8'ha3)) || ((forvar14 * reg37) != {reg24})) ?
                      {$signed(forvar13),
                          ($signed(reg34) <= $signed(reg28))} : {reg28[(4'h8):(4'h8)]}));
              reg36 <= wire0;
            end
        end
      for (forvar38 = (1'h0); (forvar38 < (1'h1)); forvar38 = (forvar38 + (1'h1)))
        begin
          for (forvar39 = (1'h0); (forvar39 < (3'h4)); forvar39 = (forvar39 + (1'h1)))
            begin
              reg40 = reg30;
              reg41 = reg20[(3'h5):(1'h1)];
              reg42 = $unsigned((reg32 + $unsigned($unsigned(((8'ha6) != reg24)))));
              reg43 <= $unsigned(reg28);
              reg44 <= reg41[(4'hb):(4'h8)];
            end
          for (forvar45 = (1'h0); (forvar45 < (3'h4)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 = $unsigned(($signed(reg27[(2'h3):(2'h2)]) ?
                  ($signed(forvar45) ?
                      (wire5 ?
                          $unsigned(wire7) : $unsigned(wire7)) : ($signed(reg28) ?
                          (reg20 ?
                              reg32 : reg15) : $unsigned(reg12))) : (&($unsigned(reg41) && $unsigned(forvar8)))));
              reg47 = (~&$signed("1xKqHy9aC"));
              reg48 <= $unsigned(reg30);
              reg49 <= ((($signed(reg17) ?
                      reg33[(4'h9):(4'h9)] : (((8'hae) != reg43) << wire0)) ?
                  (^~$unsigned(forvar8[(3'h4):(1'h0)])) : $unsigned((|reg42))) && $unsigned({((^forvar39) ?
                      {forvar19, forvar38} : $unsigned((8'h9e)))}));
            end
        end
      reg50 = $unsigned((!$unsigned(reg16[(3'h5):(2'h2)])));
    end
  module51 modinst558 (wire557, clk, reg21, reg25, forvar23, reg20);
  assign wire559 = (+reg44);
  assign wire560 = (forvar13[(2'h3):(1'h1)] ?
                       ($unsigned(reg46) ?
                           (reg21 ?
                               (wire2 ?
                                   (~|forvar23) : (wire559 ?
                                       reg49 : reg25)) : $unsigned({reg22})) : $signed((!(forvar39 ?
                               wire2 : (7'h44))))) : reg22);
  assign wire561 = reg41;
  always
    @(posedge clk) begin
      if (wire7)
        begin
          reg562 = ($unsigned(("itAVTS6Jn" <= (forvar18 <<< (&reg37)))) == (reg15[(1'h0):(1'h0)] ^~ ((~|reg37[(1'h1):(1'h0)]) ^~ ({reg30,
                  reg16} ?
              wire6 : $signed(reg50)))));
          if ($signed(forvar8[(4'hb):(3'h4)]))
            begin
              reg563 <= "";
              reg564 = {({($signed(wire559) ?
                          $unsigned((8'hb3)) : $signed(reg48))} > reg40)};
            end
          else
            begin
              reg563 <= (!(~((((8'ha4) ^~ reg42) == $unsigned(wire3)) << ($signed(reg42) || (8'hb2)))));
            end
        end
      else
        begin
          for (forvar562 = (1'h0); (forvar562 < (3'h4)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 = ((&wire557) ?
                  $signed(forvar39[(3'h4):(2'h2)]) : (8'h9c));
              reg564 <= reg33[(2'h2):(1'h1)];
            end
          for (forvar565 = (1'h0); (forvar565 < (1'h0)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg566 <= $signed($unsigned($unsigned($signed((-reg36)))));
            end
          for (forvar567 = (1'h0); (forvar567 < (3'h4)); forvar567 = (forvar567 + (1'h1)))
            begin
              reg568 = reg48[(3'h4):(1'h1)];
              reg569 <= (&$signed({(8'hb2)}));
              reg570 <= ((~&$signed(reg17[(4'ha):(3'h7)])) ~^ ((($unsigned(reg564) ?
                          wire5 : (!wire2)) ?
                      $unsigned($signed(reg48)) : (|(&reg16))) ?
                  wire3[(1'h1):(1'h0)] : ((reg25 ?
                      reg17[(3'h7):(2'h2)] : $signed(reg11)) - {forvar567,
                      ((8'ha8) ? wire5 : reg15)})));
              reg571 <= "pdlm7dTiKZqfm";
            end
          for (forvar572 = (1'h0); (forvar572 < (1'h0)); forvar572 = (forvar572 + (1'h1)))
            begin
              reg573 <= ((reg11[(3'h4):(1'h0)] <<< $unsigned(((~|forvar14) - $unsigned(forvar26)))) ?
                  forvar565 : $signed((reg571[(4'h8):(2'h3)] >> $signed(reg47[(5'h12):(3'h5)]))));
              reg574 = ({(-forvar562),
                  "CIp264caXNW71OTi"} < $signed(reg40[(3'h5):(3'h5)]));
              reg575 = forvar19[(3'h7):(3'h7)];
              reg576 = (~|($signed(reg564) ?
                  (reg47 ? reg50 : $unsigned((~wire560))) : reg573));
              reg577 <= (&forvar18);
            end
        end
      if (($unsigned("Hy5JeB7ib") ?
          ($unsigned((~|{(8'hb4), forvar18})) ?
              ($signed((reg577 ?
                  wire1 : reg564)) >> forvar14) : reg31[(2'h2):(1'h0)]) : {$unsigned(reg30)}))
        begin
          for (forvar578 = (1'h0); (forvar578 < (2'h3)); forvar578 = (forvar578 + (1'h1)))
            begin
              reg579 = $signed($unsigned((($unsigned(reg33) != (forvar572 ?
                      reg41 : wire559)) ?
                  (-((8'hae) ?
                      forvar14 : wire5)) : $signed((forvar26 | (8'ha4))))));
              reg580 = (&$unsigned(($signed(reg575) ?
                  (+(reg30 ? forvar38 : reg31)) : reg46)));
              reg581 = $signed({((~&forvar19[(4'h8):(1'h1)]) ?
                      (reg41 ?
                          reg566[(1'h0):(1'h0)] : (~|reg46)) : $unsigned($unsigned(reg580))),
                  $signed(reg562)});
              reg582 <= ({(~^reg581[(4'h8):(3'h5)]),
                  {"H7YPpOVVQ8eKUXktUB", (~&{forvar578, reg574})}} <<< (8'hb3));
            end
          reg583 = (reg49[(2'h3):(2'h2)] >= reg41[(4'hc):(3'h6)]);
          reg584 <= (+$signed(($signed($signed(reg579)) * reg36)));
        end
      else
        begin
          if ((8'hb3))
            begin
              reg578 <= (reg30[(2'h2):(1'h1)] ?
                  $unsigned(({$unsigned(forvar10)} ?
                      $signed($signed(reg25)) : $unsigned((reg580 ^~ forvar45)))) : $unsigned((forvar13 != $unsigned({reg35}))));
              reg579 = ("E" ?
                  (~{forvar26,
                      ((wire2 ? forvar45 : reg32) ?
                          (forvar26 <= reg48) : $unsigned((8'ha0)))}) : reg46);
            end
          else
            begin
              reg578 = reg44[(4'hc):(3'h7)];
              reg579 = $signed({(-(~^reg49[(1'h0):(1'h0)]))});
              reg580 <= (reg36[(2'h2):(1'h1)] >> {reg583});
              reg581 = forvar13;
            end
          for (forvar582 = (1'h0); (forvar582 < (1'h1)); forvar582 = (forvar582 + (1'h1)))
            begin
              reg583 <= {reg50[(1'h0):(1'h0)],
                  (({reg579} * $unsigned($signed(reg579))) ?
                      ((~&reg21[(4'h8):(2'h3)]) > $unsigned($signed(wire560))) : (&"ZZbwAnQ5Ku064LC2JoE"))};
              reg584 <= {reg31};
              reg585 <= ((+(($signed(reg11) ^~ wire560[(1'h0):(1'h0)]) ?
                  $unsigned(forvar13[(4'h8):(1'h1)]) : (~&$signed(forvar565)))) && wire560);
              reg586 <= ((reg573[(3'h7):(3'h4)] ?
                      wire559 : ($signed(forvar23[(2'h2):(1'h0)]) <= $unsigned(forvar38[(1'h1):(1'h1)]))) ?
                  reg580 : $signed(reg566));
            end
        end
      reg587 = (8'h9c);
      for (forvar588 = (1'h0); (forvar588 < (2'h2)); forvar588 = (forvar588 + (1'h1)))
        begin
          if (((+$unsigned(($unsigned(reg580) <<< (reg22 ?
                  wire559 : (8'hb7))))) ?
              forvar18 : (^reg44)))
            begin
              reg589 = (8'hb2);
              reg590 = "pa61rGl";
              reg591 <= $unsigned(wire1);
            end
          else
            begin
              reg589 <= reg34;
              reg590 <= reg17[(5'h10):(2'h2)];
              reg591 <= {$signed((~$unsigned({forvar45})))};
            end
          for (forvar592 = (1'h0); (forvar592 < (1'h1)); forvar592 = (forvar592 + (1'h1)))
            begin
              reg593 = forvar578;
              reg594 <= forvar19[(2'h3):(2'h2)];
            end
          for (forvar595 = (1'h0); (forvar595 < (3'h4)); forvar595 = (forvar595 + (1'h1)))
            begin
              reg596 = ((((reg578 ?
                  $signed((8'ha5)) : $signed((8'h9c))) != {(reg40 ?
                      (8'ha7) : reg590),
                  {reg47, (7'h40)}}) + ($unsigned((-wire3)) ?
                  ("Wl" ?
                      $unsigned(reg29) : reg585[(1'h1):(1'h1)]) : {$signed(forvar13)})) ~^ reg579[(3'h7):(2'h3)]);
              reg597 = $signed($unsigned((^~$signed(reg16[(1'h1):(1'h0)]))));
              reg598 = reg11;
              reg599 <= ((8'haa) ?
                  reg582 : (&$unsigned((reg48[(2'h3):(2'h3)] ?
                      (reg586 > reg596) : (8'hbc)))));
              reg600 = forvar582[(4'h9):(4'h9)];
            end
          reg601 <= $unsigned((8'hb7));
        end
      for (forvar602 = (1'h0); (forvar602 < (3'h4)); forvar602 = (forvar602 + (1'h1)))
        begin
          for (forvar603 = (1'h0); (forvar603 < (1'h0)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= (8'hb9);
              reg605 <= $unsigned($signed(((~^"qdmfRDqrUup02Yfpi") + (8'hb7))));
              reg606 = (7'h40);
              reg607 = $unsigned((~&forvar39[(3'h4):(2'h3)]));
            end
          for (forvar608 = (1'h0); (forvar608 < (1'h1)); forvar608 = (forvar608 + (1'h1)))
            begin
              reg609 <= ((((|reg571) ~^ "P51OXUxnuLuV9A1") ?
                      reg34[(4'h8):(3'h7)] : $unsigned(reg48)) ?
                  reg35[(4'hd):(4'ha)] : ($unsigned(({wire6,
                          reg584} && reg584[(4'h8):(3'h5)])) ?
                      $unsigned((reg46[(4'hf):(4'ha)] ?
                          {reg43} : reg569[(3'h4):(1'h0)])) : (~&forvar45[(3'h5):(2'h2)])));
            end
          reg610 = reg42[(5'h15):(3'h4)];
          for (forvar611 = (1'h0); (forvar611 < (3'h4)); forvar611 = (forvar611 + (1'h1)))
            begin
              reg612 <= (($signed((^~$unsigned(reg589))) ~^ (reg562[(3'h5):(1'h1)] ?
                  reg610 : reg571[(4'he):(3'h5)])) <<< reg563[(3'h4):(1'h0)]);
              reg613 <= $unsigned({(($signed(forvar565) ?
                      $unsigned(forvar578) : (reg20 ?
                          wire557 : forvar14)) << $signed((forvar602 ?
                      reg587 : reg34))),
                  $unsigned(((reg586 ^ (8'hae)) ? wire0 : $signed(reg607)))});
              reg614 = $signed($unsigned({((&wire559) != $signed((8'ha6))),
                  ($unsigned(reg587) || {reg40, reg571})}));
            end
        end
    end
  module615 modinst843 (.y(wire842), .wire618(wire7), .clk(clk), .wire616(forvar8), .wire619(forvar45), .wire617(reg17), .wire620(wire559));
  always
    @(posedge clk) begin
      reg844 <= (8'hb6);
      if (($signed(forvar611[(3'h4):(2'h3)]) ?
          ($signed(reg613) | (8'hb3)) : "svI3i9Gq9UO9RDYE"))
        begin
          reg845 <= $unsigned(forvar19);
          for (forvar846 = (1'h0); (forvar846 < (2'h3)); forvar846 = (forvar846 + (1'h1)))
            begin
              reg847 = $unsigned((reg16 > reg590[(2'h3):(2'h2)]));
              reg848 = (^~"svnl");
              reg849 = forvar23;
            end
          reg850 = ((8'hbf) ~^ $signed(forvar45[(1'h0):(1'h0)]));
          reg851 = $unsigned(forvar592[(5'h15):(5'h12)]);
          for (forvar852 = (1'h0); (forvar852 < (1'h0)); forvar852 = (forvar852 + (1'h1)))
            begin
              reg853 <= $signed(($unsigned((~^forvar23[(3'h7):(3'h7)])) ?
                  ($unsigned($signed(wire557)) <= ($unsigned(forvar19) ?
                      (reg581 ?
                          forvar45 : reg46) : (8'hb4))) : reg600[(2'h2):(1'h0)]));
              reg854 = {$signed($unsigned(reg583))};
              reg855 = ($signed($unsigned($unsigned(reg36[(2'h3):(1'h0)]))) ?
                  {((~reg594) ? "" : "mGwN")} : reg610);
              reg856 <= reg586;
              reg857 = $unsigned((~^$signed(reg16[(3'h5):(1'h1)])));
            end
        end
      else
        begin
          for (forvar845 = (1'h0); (forvar845 < (1'h1)); forvar845 = (forvar845 + (1'h1)))
            begin
              reg846 = ($unsigned(("Rcu6wf20ra8Hg" ~^ $unsigned((reg564 ?
                      (8'h9e) : reg599)))) ?
                  $signed($unsigned($unsigned(forvar14))) : $unsigned("K7"));
              reg847 <= reg12[(3'h6):(3'h4)];
              reg848 = (~|{{(|((8'ha5) >> forvar38))}});
              reg849 = reg856[(3'h7):(1'h1)];
              reg850 = forvar45[(2'h2):(1'h0)];
            end
          for (forvar851 = (1'h0); (forvar851 < (2'h2)); forvar851 = (forvar851 + (1'h1)))
            begin
              reg852 = (^($signed(reg12) ?
                  {(reg12 ? $unsigned(reg573) : $unsigned((7'h41))),
                      (reg15 ? (+forvar852) : (8'ha3))} : ({((8'h9f) ?
                              reg576 : forvar18),
                          $unsigned(reg586)} ?
                      forvar565[(2'h2):(1'h1)] : wire1[(3'h4):(1'h1)])));
              reg853 = $unsigned($signed(reg569));
              reg854 = $unsigned($signed(reg610));
              reg855 = ({reg576, forvar588[(3'h6):(3'h5)]} + (|({reg46} ?
                  (^~$unsigned(reg577)) : forvar608)));
            end
        end
      for (forvar858 = (1'h0); (forvar858 < (1'h0)); forvar858 = (forvar858 + (1'h1)))
        begin
          reg859 = {$unsigned($unsigned(reg12)),
              (forvar39[(4'h8):(4'h8)] ?
                  forvar578[(4'h8):(3'h5)] : $unsigned((((8'hbd) && (7'h41)) <<< (~|reg845))))};
          for (forvar860 = (1'h0); (forvar860 < (1'h0)); forvar860 = (forvar860 + (1'h1)))
            begin
              reg861 <= {($signed(reg16) | wire557)};
              reg862 = (+forvar10[(2'h2):(2'h2)]);
              reg863 <= (7'h43);
            end
          reg864 <= wire559[(5'h10):(2'h2)];
        end
      reg865 <= (($unsigned(reg12) >>> (((forvar608 ? forvar567 : wire1) ?
              wire5 : reg35[(4'hf):(4'he)]) ?
          ((reg846 | reg852) ?
              $unsigned(reg563) : forvar602[(2'h3):(1'h1)]) : $unsigned($signed(reg21)))) || $signed({forvar19[(4'hd):(3'h6)]}));
    end
  always
    @(posedge clk) begin
      for (forvar866 = (1'h0); (forvar866 < (1'h1)); forvar866 = (forvar866 + (1'h1)))
        begin
          for (forvar867 = (1'h0); (forvar867 < (1'h0)); forvar867 = (forvar867 + (1'h1)))
            begin
              reg868 = $signed($unsigned($unsigned((~&$signed(reg574)))));
            end
          for (forvar869 = (1'h0); (forvar869 < (1'h1)); forvar869 = (forvar869 + (1'h1)))
            begin
              reg870 = reg35[(3'h4):(2'h3)];
              reg871 <= ((8'hb9) - $unsigned(({(reg845 * forvar852),
                  (reg856 ? reg48 : forvar572)} | ("sUInEHursd4vqd" ?
                  reg850[(4'hb):(3'h5)] : (reg613 ? reg564 : forvar578)))));
              reg872 <= $unsigned((((&{reg32}) && (reg593 ?
                      $unsigned((7'h43)) : (reg593 ^ forvar18))) ?
                  forvar26[(3'h6):(2'h3)] : ((8'ha3) - reg24)));
              reg873 = $unsigned((-reg598));
            end
          for (forvar874 = (1'h0); (forvar874 < (2'h2)); forvar874 = (forvar874 + (1'h1)))
            begin
              reg875 = reg30[(2'h2):(1'h0)];
              reg876 <= (reg875[(4'hd):(4'hc)] ?
                  (($signed(reg586) ?
                      reg601 : "YnY4WYUrAP6Lk3pGpsHl") ^ (reg605[(3'h4):(2'h2)] ?
                      forvar23[(3'h7):(3'h4)] : (&((7'h44) ?
                          reg609 : reg598)))) : {(8'h9e),
                      $signed(((forvar608 ? reg574 : forvar603) <= (wire557 ?
                          reg582 : reg25)))});
            end
          if ((reg29 ?
              ((($unsigned(reg581) || (~reg605)) == reg855[(3'h4):(1'h0)]) == $unsigned((8'ha5))) : $signed((!((&forvar8) ?
                  forvar845 : $signed(reg599))))))
            begin
              reg877 <= ((reg609 >= {$unsigned(reg871[(4'ha):(3'h7)])}) >> (~&$unsigned($signed({reg40,
                  reg21}))));
              reg878 = (~|(+(~$unsigned((reg28 ? reg50 : (8'hb4))))));
            end
          else
            begin
              reg877 = {(8'ha4)};
              reg878 <= ($unsigned($signed($signed({forvar23, reg46}))) ?
                  (reg851[(1'h1):(1'h1)] ?
                      reg24[(4'ha):(3'h5)] : ((+$unsigned((8'hbe))) << $signed($signed((8'hb5))))) : $signed(reg581));
            end
        end
      for (forvar879 = (1'h0); (forvar879 < (1'h1)); forvar879 = (forvar879 + (1'h1)))
        begin
          reg880 = reg848[(4'h9):(3'h6)];
        end
    end
  always
    @(posedge clk) begin
      reg881 <= {wire5};
    end
  module708 modinst883 (wire882, clk, forvar45, forvar23, wire560, reg600, forvar852);
  always
    @(posedge clk) begin
      for (forvar884 = (1'h0); (forvar884 < (1'h1)); forvar884 = (forvar884 + (1'h1)))
        begin
          reg885 = reg28;
          for (forvar886 = (1'h0); (forvar886 < (3'h4)); forvar886 = (forvar886 + (1'h1)))
            begin
              reg887 <= wire7;
              reg888 = forvar588[(3'h7):(3'h6)];
              reg889 <= (~&((-{reg852[(2'h3):(2'h2)],
                  {reg871, reg22}}) > ((-reg607) && {(!reg22),
                  $unsigned((8'haa))})));
              reg890 <= reg872[(4'ha):(3'h7)];
              reg891 <= (((($unsigned(wire557) ?
                  reg47 : {reg872,
                      reg606}) - (reg562[(3'h6):(1'h0)] & (+reg877))) - reg580) & forvar567[(5'h14):(5'h10)]);
            end
          for (forvar892 = (1'h0); (forvar892 < (1'h1)); forvar892 = (forvar892 + (1'h1)))
            begin
              reg893 = (8'haa);
              reg894 <= (($unsigned((-$unsigned(reg42))) >= (|$unsigned({reg872}))) ?
                  (~^wire2) : $unsigned((+$signed($unsigned(reg580)))));
              reg895 = $unsigned({(&reg612)});
              reg896 = ($signed($signed($signed($unsigned(reg890)))) ?
                  (reg610[(3'h7):(3'h7)] ?
                      {($signed((8'ha1)) ?
                              (wire3 <<< (8'hbf)) : $signed(reg597))} : reg574[(4'hb):(4'ha)]) : reg601);
              reg897 = $signed({(&forvar602[(3'h4):(1'h1)]), (!(|(&reg42)))});
            end
        end
      reg898 = $signed(($signed((reg609 ?
              {wire3, forvar860} : $unsigned(wire1))) ?
          reg577 : $signed(((8'ha1) < wire6[(3'h6):(3'h4)]))));
      for (forvar899 = (1'h0); (forvar899 < (1'h1)); forvar899 = (forvar899 + (1'h1)))
        begin
          for (forvar900 = (1'h0); (forvar900 < (2'h3)); forvar900 = (forvar900 + (1'h1)))
            begin
              reg901 = (reg852[(3'h6):(2'h3)] || (~^forvar38[(3'h5):(2'h3)]));
              reg902 = $unsigned(($unsigned((wire557[(4'hb):(1'h1)] ?
                      (forvar595 || forvar900) : $unsigned(reg590))) ?
                  (^(reg844[(2'h2):(1'h1)] && (!forvar14))) : (($signed(reg851) ?
                      $signed(wire842) : $unsigned(reg16)) > {$unsigned(forvar869)})));
              reg903 <= reg41;
            end
          for (forvar904 = (1'h0); (forvar904 < (1'h0)); forvar904 = (forvar904 + (1'h1)))
            begin
              reg905 = (forvar879[(4'he):(1'h0)] ?
                  (($unsigned((reg566 ? (8'ha4) : (8'ha1))) ?
                      $signed((!reg901)) : ((reg37 ? (8'h9e) : wire2) ?
                          {forvar879,
                              reg845} : reg589)) == ((!$signed(forvar851)) ?
                      (forvar565[(4'hd):(2'h2)] == "No5m3YcPir7Mi1VFzT") : $unsigned(reg50[(1'h1):(1'h1)]))) : forvar603[(4'hd):(3'h4)]);
              reg906 <= {$signed((!reg569[(1'h1):(1'h1)]))};
            end
          reg907 <= forvar38;
        end
    end
  assign wire908 = wire3[(4'hd):(4'hd)];
  assign wire909 = (^(|(&reg848)));
  assign wire910 = $unsigned(forvar565[(3'h6):(2'h2)]);
  assign wire911 = $unsigned(reg845);
  module326 modinst913 (.wire329(reg891), .wire331(reg600), .clk(clk), .wire328(reg854), .wire330(reg889), .wire327(reg902), .y(wire912));
  always
    @(posedge clk) begin
      for (forvar914 = (1'h0); (forvar914 < (2'h3)); forvar914 = (forvar914 + (1'h1)))
        begin
          if ($unsigned($unsigned($unsigned($unsigned((reg891 ?
              reg581 : reg29))))))
            begin
              reg915 <= (((-$unsigned((|wire842))) ?
                  $unsigned(reg36[(5'h10):(3'h4)]) : (((wire911 >> (8'ha9)) ?
                      reg604[(1'h0):(1'h0)] : $signed(reg35)) ~^ $unsigned(reg601[(1'h0):(1'h0)]))) ^~ reg902);
              reg916 <= forvar578;
              reg917 <= $unsigned(((($unsigned(reg562) ^~ {reg50, reg885}) ?
                  reg872[(2'h3):(1'h1)] : wire7[(3'h6):(2'h3)]) ~^ (((7'h40) >= $unsigned((8'hbc))) && $signed("nN8PHfndd"))));
              reg918 <= reg581;
            end
          else
            begin
              reg915 = wire2[(4'hb):(4'h9)];
            end
        end
      if (($unsigned(reg890[(1'h0):(1'h0)]) ?
          $unsigned({($signed(forvar562) < "u8gPQa"),
              $signed($signed(reg15))}) : (~^(reg48[(3'h4):(1'h1)] ?
              (~&$signed(forvar13)) : $unsigned((reg850 ?
                  (8'ha0) : wire559))))))
        begin
          for (forvar919 = (1'h0); (forvar919 < (2'h3)); forvar919 = (forvar919 + (1'h1)))
            begin
              reg920 <= (reg576[(4'hf):(4'he)] ?
                  wire3[(5'h12):(3'h5)] : $unsigned((($unsigned(reg849) ?
                          (|reg613) : $signed(forvar608)) ?
                      {(reg876 ? reg583 : reg861)} : reg893)));
              reg921 <= (-("bzEo6FdBK" ?
                  ("OS42deTo0R7Ad1ed" <<< reg850[(4'hf):(4'hf)]) : (-$unsigned($unsigned(reg584)))));
              reg922 = $signed($signed((~^$signed((reg851 ?
                  (8'hb2) : (8'hb7))))));
              reg923 = reg871;
              reg924 = {(reg856[(3'h6):(3'h5)] <<< $unsigned(forvar904[(4'h8):(1'h0)]))};
            end
          for (forvar925 = (1'h0); (forvar925 < (2'h3)); forvar925 = (forvar925 + (1'h1)))
            begin
              reg926 = $signed((~"KJbGo1w"));
              reg927 <= ((|reg48[(1'h0):(1'h0)]) >>> (reg888[(1'h0):(1'h0)] || $unsigned($unsigned((reg609 ?
                  forvar851 : wire910)))));
              reg928 = reg889[(2'h3):(2'h3)];
            end
          reg929 = ($unsigned((reg48 || reg903[(4'h8):(1'h0)])) ?
              $unsigned($signed((~|$unsigned(reg614)))) : ({reg596[(4'h8):(3'h4)]} <<< reg921));
          for (forvar930 = (1'h0); (forvar930 < (3'h4)); forvar930 = (forvar930 + (1'h1)))
            begin
              reg931 <= (reg864[(4'hf):(4'hd)] > ("qf" >>> (^(reg573 ?
                  reg857[(2'h3):(2'h2)] : "q3eLrCr"))));
              reg932 = $signed(reg604[(1'h1):(1'h0)]);
              reg933 <= reg584[(4'ha):(1'h1)];
            end
          for (forvar934 = (1'h0); (forvar934 < (1'h0)); forvar934 = (forvar934 + (1'h1)))
            begin
              reg935 <= ($signed({reg873[(1'h1):(1'h1)],
                  {(reg875 ? reg898 : wire557),
                      (forvar925 ? (7'h40) : reg562)}}) > $signed(((^~(reg926 ?
                  reg609 : forvar930)) + ($unsigned(reg916) > $signed(reg931)))));
              reg936 = (~&(wire0 ?
                  $signed(((&wire909) != (~|forvar611))) : reg585[(3'h6):(2'h3)]));
            end
        end
      else
        begin
          if (forvar14)
            begin
              reg919 <= (forvar10 ?
                  (^$unsigned($unsigned("o9diLKs3KzMLPk"))) : reg876[(3'h4):(2'h2)]);
              reg920 = reg17[(4'he):(4'hb)];
              reg921 <= (~&$unsigned({(8'hae), $signed($signed(wire910))}));
              reg922 = reg919;
            end
          else
            begin
              reg919 <= reg896;
            end
          for (forvar923 = (1'h0); (forvar923 < (1'h1)); forvar923 = (forvar923 + (1'h1)))
            begin
              reg924 <= $signed(reg21);
              reg925 = forvar13;
            end
          if ($signed($signed(("9L7" ? (^~reg49) : reg848[(4'h9):(1'h0)]))))
            begin
              reg926 = $unsigned($signed((reg855 ?
                  forvar930[(2'h3):(2'h3)] : $signed({forvar10, reg889}))));
              reg927 <= $signed(("sfHOocz9TM" ?
                  (+reg610[(4'h9):(1'h0)]) : (+$signed($signed(reg566)))));
              reg928 <= forvar852[(3'h7):(2'h2)];
              reg929 = reg852[(3'h6):(2'h3)];
            end
          else
            begin
              reg926 = ({reg613[(1'h0):(1'h0)],
                      ($unsigned(forvar595) ?
                          ((reg845 <= (8'hb2)) ?
                              (reg907 ?
                                  reg931 : (8'ha2)) : (~&reg571)) : $signed((7'h42)))} ?
                  ((reg920 < reg564[(3'h4):(2'h2)]) ?
                      ((-{reg586}) << (!(reg872 && reg875))) : "Gg7qi3aqXenA28D") : {(reg33 ?
                          $unsigned($signed((8'ha4))) : $signed((|forvar884)))});
              reg927 <= $signed((((reg868[(2'h2):(1'h0)] ^ reg569) ?
                  (&(8'h9e)) : reg865[(3'h4):(2'h2)]) | "Kn8r0"));
              reg928 <= $unsigned(forvar10[(2'h3):(1'h0)]);
              reg929 <= {(wire3 ? reg579 : (8'hb5))};
            end
        end
      for (forvar937 = (1'h0); (forvar937 < (2'h3)); forvar937 = (forvar937 + (1'h1)))
        begin
          if ($unsigned($signed((-wire910[(1'h1):(1'h0)]))))
            begin
              reg938 <= $signed({(reg845 ^~ ($unsigned((7'h44)) ?
                      wire6 : wire560))});
              reg939 <= $signed($signed($unsigned($signed(reg569))));
              reg940 <= (~^($unsigned(reg587[(4'h9):(4'h8)]) + (8'hb8)));
              reg941 <= (reg600 ?
                  $unsigned($unsigned((|(reg610 ?
                      (8'h9e) : (8'hbf))))) : $signed(({$signed(forvar904),
                          {(7'h44)}} ?
                      $signed(((8'haa) ?
                          reg587 : reg844)) : $unsigned(reg601))));
              reg942 = reg918[(2'h2):(2'h2)];
            end
          else
            begin
              reg938 <= ((forvar562[(2'h3):(1'h0)] <<< reg889) ?
                  $unsigned(reg929) : (reg35 < (8'hbf)));
              reg939 = ({reg21} ?
                  ($signed(((~forvar860) ?
                      $unsigned((8'hb3)) : reg35)) <= $unsigned((&"mRZh"))) : {(8'hb6),
                      ($unsigned(forvar866) ?
                          $unsigned(reg570[(2'h2):(2'h2)]) : reg844[(2'h2):(1'h1)])});
              reg940 <= ($unsigned({$signed((forvar899 ^~ wire559))}) ?
                  {{$signed((forvar588 * forvar8))}} : (8'ha2));
              reg941 <= $unsigned(forvar884);
            end
        end
      for (forvar943 = (1'h0); (forvar943 < (1'h0)); forvar943 = (forvar943 + (1'h1)))
        begin
          for (forvar944 = (1'h0); (forvar944 < (1'h1)); forvar944 = (forvar944 + (1'h1)))
            begin
              reg945 = $signed((+($signed($signed(forvar874)) < $signed(wire908))));
              reg946 <= (^"");
              reg947 <= ($unsigned(($signed(reg597) > reg887)) >>> reg864[(4'he):(2'h2)]);
              reg948 <= $unsigned((^{(reg574 ^ (reg922 ? reg42 : reg584))}));
            end
          if ({(&((reg922 ? forvar8[(5'h11):(3'h4)] : (^~reg21)) ?
                  $unsigned((reg35 != (8'hb4))) : ($unsigned((7'h42)) ~^ (reg942 ?
                      (8'hb2) : reg921)))),
              "LmCsEvPgq6rbUY"})
            begin
              reg949 = reg563[(2'h2):(2'h2)];
              reg950 <= $unsigned((&$unsigned((forvar608[(5'h14):(4'hf)] ^~ (reg568 ?
                  reg919 : (8'ha6))))));
              reg951 <= {((-reg933) ?
                      ((-((8'hb0) < reg936)) > $signed(forvar23)) : ((reg928[(3'h4):(3'h4)] * reg42) < reg34[(1'h1):(1'h0)])),
                  "t45nkU3xS4yelx"};
              reg952 <= (((reg609[(2'h2):(2'h2)] ?
                          $signed(reg589[(1'h1):(1'h0)]) : reg852) ?
                      reg590 : (reg846[(2'h2):(1'h1)] >>> $unsigned((-forvar18)))) ?
                  (~$unsigned((^~(reg935 <= (7'h41))))) : $unsigned((~&($signed(reg923) + (reg875 ?
                      (8'hab) : (8'hb4))))));
              reg953 <= reg597[(4'hf):(3'h4)];
            end
          else
            begin
              reg949 = (|$unsigned($unsigned(forvar858[(1'h0):(1'h0)])));
              reg950 = wire912;
            end
          reg954 <= (~{("w6vgmRwB6hYK" | $unsigned($unsigned(reg895))),
              reg48[(3'h4):(2'h3)]});
          for (forvar955 = (1'h0); (forvar955 < (2'h3)); forvar955 = (forvar955 + (1'h1)))
            begin
              reg956 = ($unsigned(((reg922[(3'h6):(1'h1)] ?
                      (reg921 ? forvar578 : reg942) : forvar852) ?
                  (((8'hbf) ? reg32 : wire911) >>> $signed((7'h42))) : {reg888,
                      {reg917, (8'hbc)}})) >> ($signed((&(-reg888))) ?
                  (^~$signed($signed(reg933))) : $unsigned($unsigned((8'hb0)))));
              reg957 <= reg564;
              reg958 = "YJYN1bTVsK5xJPB0GK";
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module615
#( parameter param841 = ((~(~|(~&{(8'hab), (8'ha5)}))) ? (8'haf) : (~^(((8'h9d) ^ ((7'h40) <<< (8'hb4))) ? {(^~(8'ha0)), ((8'haa) > (8'ha7))} : {((8'ha5) || (8'had))}))) )
(y, clk, wire616, wire617, wire618, wire619, wire620);
  output wire [(32'h508):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire616;
  input wire signed [(4'hf):(1'h0)] wire617;
  input wire [(3'h7):(1'h0)] wire618;
  input wire signed [(3'h6):(1'h0)] wire619;
  input wire [(5'h14):(1'h0)] wire620;
  reg signed [(2'h2):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar837 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg836 = (1'h0);
  reg [(2'h2):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar833 = (1'h0);
  reg [(3'h7):(1'h0)] reg834 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg833 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg832 = (1'h0);
  reg [(5'h15):(1'h0)] reg831 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg830 = (1'h0);
  reg [(2'h3):(1'h0)] reg829 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg828 = (1'h0);
  reg [(4'hd):(1'h0)] reg827 = (1'h0);
  reg [(4'hc):(1'h0)] reg826 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg825 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg824 = (1'h0);
  reg [(5'h10):(1'h0)] forvar823 = (1'h0);
  reg [(5'h11):(1'h0)] reg822 = (1'h0);
  reg [(5'h15):(1'h0)] reg821 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar820 = (1'h0);
  reg [(4'he):(1'h0)] forvar819 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg818 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg817 = (1'h0);
  reg [(2'h2):(1'h0)] reg816 = (1'h0);
  reg [(2'h2):(1'h0)] reg815 = (1'h0);
  reg [(5'h14):(1'h0)] forvar814 = (1'h0);
  reg [(2'h3):(1'h0)] reg813 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire812;
  wire [(4'he):(1'h0)] wire811;
  wire [(5'h14):(1'h0)] wire621;
  reg [(4'hb):(1'h0)] forvar622 = (1'h0);
  reg [(4'hf):(1'h0)] reg623 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar624 = (1'h0);
  reg [(3'h5):(1'h0)] reg625 = (1'h0);
  reg signed [(4'he):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg628 = (1'h0);
  reg [(3'h7):(1'h0)] reg629 = (1'h0);
  reg [(3'h4):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar631 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg632 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg633 = (1'h0);
  reg [(2'h2):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg635 = (1'h0);
  reg [(4'hb):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg637 = (1'h0);
  reg [(2'h3):(1'h0)] reg638 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg639 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar640 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg642 = (1'h0);
  reg [(5'h10):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg644 = (1'h0);
  reg [(2'h3):(1'h0)] reg645 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar646 = (1'h0);
  reg [(4'hb):(1'h0)] reg647 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg648 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg649 = (1'h0);
  reg [(4'ha):(1'h0)] reg646 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg650 = (1'h0);
  reg [(4'h8):(1'h0)] reg651 = (1'h0);
  reg [(2'h2):(1'h0)] reg652 = (1'h0);
  reg [(5'h14):(1'h0)] forvar653 = (1'h0);
  reg [(5'h11):(1'h0)] reg654 = (1'h0);
  reg [(4'hd):(1'h0)] reg655 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg656 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar657 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar658 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg659 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg660 = (1'h0);
  reg [(3'h6):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar662 = (1'h0);
  reg [(2'h2):(1'h0)] reg663 = (1'h0);
  reg [(4'ha):(1'h0)] reg664 = (1'h0);
  reg signed [(4'he):(1'h0)] reg665 = (1'h0);
  reg [(5'h15):(1'h0)] forvar666 = (1'h0);
  reg signed [(4'he):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg669 = (1'h0);
  reg [(4'h9):(1'h0)] forvar670 = (1'h0);
  reg [(2'h2):(1'h0)] forvar671 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg673 = (1'h0);
  reg [(3'h4):(1'h0)] reg674 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg675 = (1'h0);
  reg [(4'h8):(1'h0)] reg676 = (1'h0);
  reg [(4'hc):(1'h0)] reg677 = (1'h0);
  reg [(3'h7):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg679 = (1'h0);
  reg [(3'h7):(1'h0)] forvar680 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg681 = (1'h0);
  reg [(4'h9):(1'h0)] reg682 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg683 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg684 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar684 = (1'h0);
  reg [(5'h10):(1'h0)] reg685 = (1'h0);
  reg [(4'hc):(1'h0)] reg686 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg687 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg689 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar690 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar691 = (1'h0);
  reg [(4'hd):(1'h0)] reg692 = (1'h0);
  reg [(3'h4):(1'h0)] reg693 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar695 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg696 = (1'h0);
  reg signed [(4'he):(1'h0)] reg697 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg698 = (1'h0);
  reg [(4'h8):(1'h0)] reg699 = (1'h0);
  reg [(3'h7):(1'h0)] reg700 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar701 = (1'h0);
  reg [(2'h2):(1'h0)] reg702 = (1'h0);
  reg [(4'hf):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg705 = (1'h0);
  reg [(4'hb):(1'h0)] reg706 = (1'h0);
  reg [(3'h4):(1'h0)] reg707 = (1'h0);
  wire [(3'h7):(1'h0)] wire809;
  assign y = {reg840,
                 reg839,
                 reg838,
                 forvar837,
                 reg836,
                 reg835,
                 forvar833,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 forvar823,
                 reg822,
                 reg821,
                 forvar820,
                 forvar819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 forvar814,
                 reg813,
                 wire812,
                 wire811,
                 wire621,
                 forvar622,
                 reg623,
                 forvar624,
                 reg625,
                 reg626,
                 reg627,
                 reg628,
                 reg629,
                 reg630,
                 forvar631,
                 reg632,
                 reg633,
                 reg634,
                 reg635,
                 reg636,
                 reg637,
                 reg638,
                 reg639,
                 forvar640,
                 reg641,
                 reg642,
                 reg643,
                 reg644,
                 reg645,
                 forvar646,
                 reg647,
                 reg648,
                 reg649,
                 reg646,
                 reg650,
                 reg651,
                 reg652,
                 forvar653,
                 reg654,
                 reg655,
                 reg656,
                 forvar657,
                 forvar658,
                 reg659,
                 reg660,
                 reg661,
                 forvar662,
                 reg663,
                 reg664,
                 reg665,
                 forvar666,
                 reg667,
                 reg668,
                 reg669,
                 forvar670,
                 forvar671,
                 reg672,
                 reg673,
                 reg674,
                 reg675,
                 reg676,
                 reg677,
                 reg678,
                 reg679,
                 forvar680,
                 reg681,
                 reg682,
                 reg683,
                 reg684,
                 forvar684,
                 reg685,
                 reg686,
                 reg687,
                 reg688,
                 reg689,
                 forvar690,
                 forvar691,
                 reg692,
                 reg693,
                 reg694,
                 forvar695,
                 reg696,
                 reg697,
                 reg698,
                 reg699,
                 reg700,
                 forvar701,
                 reg702,
                 reg703,
                 reg704,
                 reg705,
                 reg706,
                 reg707,
                 wire809,
                 (1'h0)};
  assign wire621 = ((wire618[(2'h2):(2'h2)] ~^ $unsigned(wire618[(1'h1):(1'h0)])) - $signed(((8'ha0) >> wire616)));
  always
    @(posedge clk) begin
      for (forvar622 = (1'h0); (forvar622 < (1'h0)); forvar622 = (forvar622 + (1'h1)))
        begin
          reg623 <= (($unsigned($signed((wire618 | forvar622))) ?
                  $unsigned(((wire621 + wire619) ^~ $unsigned(wire620))) : wire616) ?
              $unsigned(($signed($signed(wire617)) || (forvar622[(4'h9):(4'h9)] ?
                  wire618[(3'h7):(3'h4)] : (wire621 | wire621)))) : ($unsigned((!$unsigned((8'ha8)))) + (((~forvar622) >> $unsigned((8'hb8))) << $signed($signed(wire616)))));
          for (forvar624 = (1'h0); (forvar624 < (2'h3)); forvar624 = (forvar624 + (1'h1)))
            begin
              reg625 = $signed({$signed(wire619),
                  (wire616[(1'h1):(1'h1)] ?
                      $signed((wire619 ?
                          forvar622 : wire621)) : (&reg623[(1'h0):(1'h0)]))});
              reg626 = $signed($unsigned(reg625[(3'h5):(2'h2)]));
              reg627 = $signed((8'h9e));
              reg628 <= $signed(($unsigned(reg625[(2'h3):(2'h3)]) ?
                  (~($unsigned(wire619) ^~ $signed(wire617))) : $signed(($signed(reg623) == wire616[(2'h3):(2'h3)]))));
              reg629 <= wire617[(3'h7):(2'h2)];
            end
          reg630 <= reg627[(4'h8):(2'h2)];
          for (forvar631 = (1'h0); (forvar631 < (1'h1)); forvar631 = (forvar631 + (1'h1)))
            begin
              reg632 = wire617;
            end
          reg633 <= $unsigned((+{$signed((reg630 ? forvar624 : reg623))}));
        end
      if ($signed(($signed(({(8'hb3), wire617} ?
          {reg625, wire616} : {forvar622})) && {wire621[(5'h14):(5'h14)],
          ($unsigned(wire617) ? (forvar624 > reg625) : $signed(wire621))})))
        begin
          reg634 = wire617[(4'hb):(3'h6)];
          reg635 = ($signed(forvar622[(2'h2):(2'h2)]) << $unsigned(reg630[(3'h4):(1'h0)]));
          reg636 <= reg625;
        end
      else
        begin
          reg634 <= $signed($unsigned($unsigned(($signed((8'hab)) ?
              ((8'h9d) ^~ (8'ha8)) : (forvar624 > reg633)))));
          if ($signed(reg630))
            begin
              reg635 = $unsigned(reg634[(2'h2):(2'h2)]);
              reg636 <= ($signed((~^((reg627 != (7'h44)) ?
                      (~&reg633) : reg630[(1'h0):(1'h0)]))) ?
                  reg634[(1'h1):(1'h0)] : (wire616 || $unsigned(forvar624)));
              reg637 = (~(reg627[(5'h11):(4'he)] | ({(reg628 == (8'ha3))} | (|{(8'hb8),
                  reg634}))));
              reg638 = reg630[(2'h3):(1'h0)];
              reg639 <= reg626;
            end
          else
            begin
              reg635 = $signed({$unsigned(wire617[(4'hf):(1'h0)])});
              reg636 = wire617;
              reg637 <= wire620[(2'h2):(1'h1)];
            end
        end
      if ((+reg630[(2'h3):(2'h2)]))
        begin
          for (forvar640 = (1'h0); (forvar640 < (2'h2)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 <= (reg632[(2'h2):(1'h0)] ?
                  (+{(~^(8'h9d)), {(!wire616)}}) : (+reg637));
              reg642 = $signed(wire616);
            end
          reg643 = ($unsigned($signed($signed($signed(wire618)))) ?
              ($unsigned(wire619[(1'h1):(1'h0)]) ?
                  ((^~{reg632, reg626}) ~^ (reg637[(2'h2):(1'h0)] ?
                      "6sSdtw" : $unsigned(reg642))) : ((^$signed(reg635)) != reg634)) : $signed(wire619[(1'h0):(1'h0)]));
          if ((~|(-({(wire621 & (8'h9c))} ?
              (reg638[(1'h1):(1'h0)] ^~ (reg633 ? reg633 : reg638)) : reg635))))
            begin
              reg644 = $unsigned($signed($signed(($signed((8'ha2)) ~^ $unsigned(wire618)))));
            end
          else
            begin
              reg644 = {$unsigned(reg628[(4'h9):(3'h6)])};
              reg645 <= reg635[(4'hb):(4'h9)];
            end
          for (forvar646 = (1'h0); (forvar646 < (2'h2)); forvar646 = (forvar646 + (1'h1)))
            begin
              reg647 <= ((({reg627} << {(~&reg639)}) ?
                      "o" : reg638[(2'h2):(1'h0)]) ?
                  $signed($unsigned((reg625[(3'h4):(1'h1)] ?
                      $signed(reg628) : (forvar640 > wire620)))) : {forvar622});
              reg648 = (-$signed($signed(((wire619 ^~ reg634) - $signed(reg625)))));
              reg649 <= $signed("3vROY");
            end
        end
      else
        begin
          for (forvar640 = (1'h0); (forvar640 < (2'h3)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 <= ((($signed({wire620}) * (~|(reg637 ?
                  reg649 : reg641))) && $signed(($unsigned((7'h42)) == $signed((8'h9e))))) <= (reg628 + reg626));
              reg642 <= ($unsigned("zW7V") ?
                  wire616[(3'h7):(1'h1)] : {(-reg644),
                      $signed((!reg642[(4'hb):(3'h6)]))});
            end
          if ((^((forvar622[(2'h3):(2'h2)] ?
                  "Q5012n" : ($unsigned(reg645) == $unsigned(reg643))) ?
              $unsigned($unsigned($unsigned(wire616))) : wire618[(3'h5):(3'h5)])))
            begin
              reg643 = (+$signed(reg647[(4'ha):(1'h0)]));
              reg644 = reg641;
              reg645 <= $unsigned(wire617);
              reg646 = forvar631[(3'h4):(2'h3)];
            end
          else
            begin
              reg643 = reg645;
              reg644 = $unsigned((reg628 ?
                  "vS8cBIdw" : wire617[(3'h7):(2'h2)]));
              reg645 <= (+forvar640);
            end
          if (("gYswbT5aO8gUJG6PhTr" ?
              $unsigned($unsigned($signed((~|reg627)))) : $unsigned(wire619)))
            begin
              reg647 <= reg647;
            end
          else
            begin
              reg647 <= ($unsigned(forvar631) ? $unsigned(reg635) : reg629);
              reg648 = $unsigned({(~(~|wire617[(4'hd):(4'hb)]))});
              reg649 = (reg623[(2'h3):(1'h1)] ^ (!$signed((wire618[(3'h7):(3'h7)] ^~ (~|reg645)))));
              reg650 <= $signed(wire619[(2'h2):(1'h0)]);
              reg651 = (wire618[(3'h4):(2'h3)] ?
                  wire617 : (({$signed((7'h44)), $signed((8'h9e))} ?
                      wire619[(2'h2):(1'h0)] : $unsigned($unsigned(reg647))) & $unsigned(((^~(8'ha3)) || $signed(reg648)))));
            end
          reg652 = reg648;
          for (forvar653 = (1'h0); (forvar653 < (2'h3)); forvar653 = (forvar653 + (1'h1)))
            begin
              reg654 = (!($signed(((reg637 && reg648) >> $signed(reg633))) ?
                  ({wire617} * ($unsigned(wire619) | wire620)) : ("ctmCfSeD6" ?
                      reg626[(4'h9):(2'h2)] : $signed(wire620))));
              reg655 = ($signed(($signed((|reg628)) >> "WhJFpxEZOi8ti")) >> (8'hac));
            end
        end
    end
  always
    @(posedge clk) begin
      reg656 <= ((~{((~^reg635) || $signed((8'had)))}) > forvar640[(1'h0):(1'h0)]);
      for (forvar657 = (1'h0); (forvar657 < (1'h0)); forvar657 = (forvar657 + (1'h1)))
        begin
          for (forvar658 = (1'h0); (forvar658 < (1'h0)); forvar658 = (forvar658 + (1'h1)))
            begin
              reg659 = $signed("yBS0");
              reg660 = forvar646;
            end
          reg661 = (reg649 + $signed(($unsigned((!reg637)) ^~ (((8'ha9) ?
              (8'haa) : forvar622) && (reg649 ? reg642 : (8'haa))))));
          for (forvar662 = (1'h0); (forvar662 < (2'h2)); forvar662 = (forvar662 + (1'h1)))
            begin
              reg663 = (7'h40);
              reg664 = (~|$signed({reg632[(2'h2):(2'h2)],
                  ($unsigned(reg627) ?
                      (reg636 ? reg644 : (8'hbe)) : (reg647 ?
                          (8'hb5) : reg639))}));
              reg665 <= ((reg660[(4'h9):(3'h6)] <= $unsigned(forvar646)) ?
                  wire621 : $signed((reg663 ^ forvar662)));
            end
          for (forvar666 = (1'h0); (forvar666 < (1'h1)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 <= (^(~|$unsigned((&reg632))));
              reg668 = reg652[(2'h2):(1'h0)];
              reg669 = $signed(((reg651[(1'h1):(1'h0)] ?
                      ((reg655 ?
                          reg628 : reg645) + $signed(reg668)) : ((8'ha4) >> forvar640[(4'ha):(3'h4)])) ?
                  ({(forvar624 ? reg645 : reg637)} | ($unsigned(reg639) ?
                      (reg634 ?
                          (8'ha1) : reg665) : (8'hb3))) : reg648[(3'h4):(2'h3)]));
            end
        end
      for (forvar670 = (1'h0); (forvar670 < (1'h0)); forvar670 = (forvar670 + (1'h1)))
        begin
          for (forvar671 = (1'h0); (forvar671 < (2'h3)); forvar671 = (forvar671 + (1'h1)))
            begin
              reg672 = $signed($unsigned(forvar640));
              reg673 <= (((+reg659) | ((^~$unsigned(forvar624)) != (forvar646 <<< ((7'h42) ^ forvar622)))) ?
                  $unsigned((+reg625)) : $signed($signed((reg667[(4'hd):(3'h4)] <= reg651[(3'h7):(2'h2)]))));
              reg674 <= wire619;
            end
          if (((|forvar662[(1'h1):(1'h1)]) ?
              (&(~&$signed((reg652 != (8'h9c))))) : reg669[(1'h0):(1'h0)]))
            begin
              reg675 = {$unsigned(wire617[(4'hd):(4'ha)])};
              reg676 = (($signed(forvar671) | $unsigned({(~|reg645)})) ?
                  (~$signed("KlqpQcwv")) : reg623[(4'h9):(4'h8)]);
              reg677 <= {{{(reg659 ? (~&forvar646) : reg659),
                          $signed((!reg625))}},
                  {(|"7pv")}};
              reg678 = ($unsigned({($unsigned(reg642) << (reg677 == reg642)),
                      ({(8'hb0), (7'h43)} <= (reg668 ? reg675 : reg665))}) ?
                  reg656 : {$unsigned($unsigned((forvar631 ~^ reg644)))});
              reg679 <= $unsigned((~|$unsigned(($signed(reg663) && $unsigned(reg627)))));
            end
          else
            begin
              reg675 = reg652;
              reg676 = $unsigned($unsigned($unsigned((~^(forvar658 ?
                  reg623 : forvar640)))));
              reg677 <= ("sgeZ28g1YyZVC" ?
                  $signed($unsigned("UafZJSHIaz16h")) : (forvar666 ?
                      $signed("R2q22lU3mo3a") : {forvar657,
                          ($unsigned(reg639) ?
                              (^forvar671) : reg638[(1'h0):(1'h0)])}));
            end
          for (forvar680 = (1'h0); (forvar680 < (3'h4)); forvar680 = (forvar680 + (1'h1)))
            begin
              reg681 = $unsigned($unsigned(wire620[(4'hd):(4'hd)]));
              reg682 <= $unsigned($signed(($signed($signed(reg648)) ?
                  reg647[(2'h3):(2'h2)] : {{reg630, wire621}})));
              reg683 <= {{$signed((-reg673[(2'h2):(1'h1)])),
                      (~^($unsigned(reg648) <= (~^forvar624)))},
                  ((7'h42) ? $unsigned(reg643) : forvar646)};
            end
        end
      if ((^~$unsigned((~&"SMNgZqRp0mn"))))
        begin
          reg684 <= $unsigned(("A38uETuO1GV3Adh" ?
              (reg642[(3'h4):(1'h0)] != $unsigned($unsigned(forvar670))) : "1"));
        end
      else
        begin
          for (forvar684 = (1'h0); (forvar684 < (2'h3)); forvar684 = (forvar684 + (1'h1)))
            begin
              reg685 <= ({{$signed((~^reg677))}} >>> $signed($unsigned((~reg682))));
              reg686 <= (+reg661);
              reg687 = (&wire619);
              reg688 <= (wire616 ?
                  $unsigned((-((reg651 ^~ (8'ha2)) ?
                      reg672 : forvar631))) : ((wire618[(3'h6):(1'h1)] ?
                          (~"bfvTTW3Gs1FbyyWn1Vbf") : $unsigned((+reg644))) ?
                      wire619 : reg659));
            end
          reg689 = reg681;
        end
      for (forvar690 = (1'h0); (forvar690 < (3'h4)); forvar690 = (forvar690 + (1'h1)))
        begin
          for (forvar691 = (1'h0); (forvar691 < (1'h0)); forvar691 = (forvar691 + (1'h1)))
            begin
              reg692 <= (reg646[(3'h5):(3'h5)] ?
                  (forvar631 ?
                      ({{forvar671}} >>> (8'hb9)) : reg627[(5'h12):(3'h7)]) : (-$signed($signed(reg673[(2'h2):(2'h2)]))));
              reg693 = forvar624;
              reg694 <= (!($signed((((8'ha7) | reg646) << (&reg669))) ?
                  forvar671[(1'h1):(1'h0)] : reg632[(4'ha):(4'h8)]));
            end
          for (forvar695 = (1'h0); (forvar695 < (3'h4)); forvar695 = (forvar695 + (1'h1)))
            begin
              reg696 <= $unsigned($signed(forvar691[(1'h0):(1'h0)]));
              reg697 <= reg686[(4'hc):(3'h5)];
              reg698 = ($signed(reg641) ?
                  $signed((reg679[(1'h1):(1'h0)] ?
                      $unsigned(reg674[(2'h3):(2'h3)]) : $signed((~&reg664)))) : (((-$signed((8'ha7))) >> {reg677[(2'h2):(2'h2)]}) ?
                      ($unsigned($unsigned(reg652)) && (reg650[(3'h7):(1'h1)] ?
                          ((8'hb1) >>> (8'had)) : (8'ha8))) : (forvar646[(2'h2):(1'h0)] != (|$signed(reg688)))));
              reg699 <= ($unsigned((~^(reg646 || reg668))) >> wire616[(2'h3):(2'h3)]);
              reg700 <= $signed((reg697[(4'he):(3'h4)] == (((~(8'hb7)) ?
                  $unsigned(reg687) : $unsigned(reg689)) <<< $signed((&reg664)))));
            end
          for (forvar701 = (1'h0); (forvar701 < (1'h1)); forvar701 = (forvar701 + (1'h1)))
            begin
              reg702 = $signed(forvar691[(3'h5):(3'h4)]);
              reg703 <= $signed($unsigned({(~&wire619)}));
              reg704 <= $unsigned((reg632 + reg686));
              reg705 = (reg649 ?
                  (~forvar622) : (+(reg678 ?
                      (8'hb4) : ($unsigned(reg673) ?
                          ((8'hb9) ?
                              (8'hb9) : reg637) : forvar680[(3'h4):(1'h0)]))));
            end
          reg706 = $signed((forvar671[(2'h2):(2'h2)] ?
              {reg651[(2'h2):(1'h0)]} : (~&reg650)));
          reg707 <= (&(!reg678));
        end
    end
  module708 modinst810 (.wire710(reg699), .wire713(reg679), .wire711(forvar684), .y(wire809), .clk(clk), .wire712(reg696), .wire709(reg689));
  assign wire811 = ((($signed(reg627) ?
                       wire617[(4'ha):(1'h0)] : $signed({wire618,
                           wire616})) + $unsigned($signed(reg687[(2'h2):(1'h1)]))) - reg646);
  assign wire812 = reg629;
  always
    @(posedge clk) begin
      reg813 = $unsigned(reg704[(4'hc):(4'ha)]);
      for (forvar814 = (1'h0); (forvar814 < (2'h2)); forvar814 = (forvar814 + (1'h1)))
        begin
          if (forvar670)
            begin
              reg815 = ($signed((~&((forvar670 ?
                      (8'hb1) : wire617) >> reg654[(1'h0):(1'h0)]))) ?
                  $unsigned(($unsigned((reg663 ^~ reg667)) - $signed({reg665,
                      reg663}))) : (({reg688[(1'h0):(1'h0)]} ^ $unsigned({reg813})) >= $unsigned((-reg707))));
              reg816 <= "66Cy58FV7Tdn2HR6FQm6";
            end
          else
            begin
              reg815 = reg649[(1'h1):(1'h0)];
              reg816 = ({(^~((~reg634) ? {reg679} : forvar624[(4'h9):(4'h9)])),
                  (((-forvar657) ?
                          forvar653[(3'h6):(2'h3)] : (reg696 ?
                              forvar684 : reg627)) ?
                      wire618 : ("naheLB" ^ (reg698 ?
                          reg685 : (8'h9c))))} <= ((-($unsigned(reg625) <= "T3Fs7YaB2YD7g2")) ?
                  $signed(($unsigned((8'ha5)) || (8'ha9))) : $unsigned(((^~reg678) ?
                      (forvar658 ? reg679 : reg664) : (reg623 <= forvar666)))));
              reg817 <= {($unsigned($signed(reg699)) >= {$signed(reg660[(3'h5):(3'h5)]),
                      $signed((^forvar701))}),
                  (reg699 <= ($unsigned(reg629[(2'h3):(1'h1)]) ?
                      ({reg674} <= (~reg696)) : $signed($unsigned(reg688))))};
              reg818 <= $unsigned($signed((^~{reg705[(3'h4):(2'h3)],
                  $signed(reg682)})));
            end
        end
      for (forvar819 = (1'h0); (forvar819 < (2'h2)); forvar819 = (forvar819 + (1'h1)))
        begin
          for (forvar820 = (1'h0); (forvar820 < (2'h3)); forvar820 = (forvar820 + (1'h1)))
            begin
              reg821 = {(!reg633[(1'h0):(1'h0)]), (^~reg628)};
            end
        end
      reg822 <= forvar695[(4'h8):(1'h1)];
      for (forvar823 = (1'h0); (forvar823 < (1'h0)); forvar823 = (forvar823 + (1'h1)))
        begin
          reg824 <= (~|{$unsigned($signed((~|reg623)))});
          if (reg684[(1'h1):(1'h1)])
            begin
              reg825 <= $unsigned((reg816 > $signed(reg668[(2'h3):(1'h1)])));
              reg826 = $unsigned((~$signed(reg693)));
              reg827 = wire812[(4'h8):(3'h7)];
              reg828 <= reg693;
            end
          else
            begin
              reg825 = (!$signed($signed($signed((forvar680 ?
                  (8'haf) : reg826)))));
              reg826 <= ((reg697 >= ({wire621, (reg693 | reg623)} ?
                      ((forvar695 ^~ (8'hb2)) + reg686[(4'hb):(4'hb)]) : {(reg649 >>> forvar657)})) ?
                  reg684[(1'h0):(1'h0)] : reg702[(1'h0):(1'h0)]);
            end
          if ((8'hba))
            begin
              reg829 <= $unsigned(wire809);
            end
          else
            begin
              reg829 <= "nxBYt";
              reg830 <= (reg642[(3'h6):(3'h6)] >= ($unsigned($signed($signed((8'ha2)))) ?
                  (|$signed((+forvar671))) : "I8kGmDJ9Vy7"));
              reg831 = forvar691[(1'h0):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed(($signed(reg688) & reg699[(3'h5):(3'h4)])))
        begin
          if ((^(8'h9d)))
            begin
              reg832 = reg648[(2'h2):(1'h0)];
              reg833 = $signed($signed(reg698[(3'h6):(3'h6)]));
              reg834 = reg646;
            end
          else
            begin
              reg832 = ($unsigned($unsigned(reg656[(2'h2):(1'h1)])) || reg832[(2'h2):(2'h2)]);
              reg833 = ($signed((+"bosANN2")) ?
                  $unsigned($signed((-(reg689 ?
                      reg833 : forvar662)))) : (&(~(+(reg636 <<< reg661)))));
              reg834 <= (($signed(reg647[(4'h9):(2'h2)]) || (wire619[(1'h0):(1'h0)] <<< $signed({reg677,
                  reg693}))) & (^~$unsigned((((8'hbe) ^~ forvar658) ?
                  reg707 : ((8'hb4) == (8'haa))))));
            end
        end
      else
        begin
          reg832 = (+((forvar657[(3'h4):(1'h1)] ?
              (-$unsigned(reg636)) : wire619) + ($signed((~reg821)) ~^ $unsigned($signed(reg645)))));
          for (forvar833 = (1'h0); (forvar833 < (2'h3)); forvar833 = (forvar833 + (1'h1)))
            begin
              reg834 = ("f9" ?
                  $signed({(&$unsigned(reg679)),
                      reg639[(2'h2):(1'h0)]}) : $unsigned($unsigned(((+reg694) ?
                      reg683[(2'h2):(1'h0)] : $signed(forvar622)))));
              reg835 <= ($signed($signed(reg667[(1'h0):(1'h0)])) | $signed(reg705));
              reg836 <= ($signed(reg683[(3'h4):(3'h4)]) ?
                  (wire619[(2'h3):(2'h2)] & $unsigned(reg826)) : (!reg654));
            end
          for (forvar837 = (1'h0); (forvar837 < (1'h0)); forvar837 = (forvar837 + (1'h1)))
            begin
              reg838 = {$unsigned($signed(({forvar631} ?
                      reg669 : {reg655, reg833})))};
            end
          reg839 = $unsigned((8'h9e));
          reg840 = reg698;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module51  (y, clk, wire52, wire53, wire54, wire55);
  output wire [(32'h672):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire52;
  input wire [(5'h11):(1'h0)] wire53;
  input wire [(2'h3):(1'h0)] wire54;
  input wire [(5'h11):(1'h0)] wire55;
  wire [(5'h12):(1'h0)] wire556;
  wire signed [(3'h6):(1'h0)] wire555;
  wire [(5'h15):(1'h0)] wire554;
  reg signed [(5'h11):(1'h0)] reg553 = (1'h0);
  reg [(4'he):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg550 = (1'h0);
  reg [(5'h11):(1'h0)] reg549 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar548 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg547 = (1'h0);
  reg [(4'hb):(1'h0)] reg546 = (1'h0);
  reg [(4'h8):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg544 = (1'h0);
  reg [(5'h14):(1'h0)] forvar543 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg542 = (1'h0);
  reg [(4'hd):(1'h0)] reg541 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg540 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar539 = (1'h0);
  reg [(5'h13):(1'h0)] forvar538 = (1'h0);
  reg [(3'h6):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar57 = (1'h0);
  reg [(5'h14):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg59 = (1'h0);
  reg signed [(4'he):(1'h0)] reg60 = (1'h0);
  reg [(5'h12):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg62 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar63 = (1'h0);
  reg [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg67 = (1'h0);
  reg [(5'h14):(1'h0)] forvar68 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg69 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar58 = (1'h0);
  reg [(4'ha):(1'h0)] forvar72 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar73 = (1'h0);
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg76 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg77 = (1'h0);
  reg [(5'h10):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg79 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg81 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar82 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg83 = (1'h0);
  reg [(3'h4):(1'h0)] reg84 = (1'h0);
  reg [(3'h6):(1'h0)] reg85 = (1'h0);
  reg [(5'h11):(1'h0)] reg86 = (1'h0);
  reg [(2'h2):(1'h0)] reg87 = (1'h0);
  reg [(2'h3):(1'h0)] forvar88 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg91 = (1'h0);
  reg [(3'h7):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar93 = (1'h0);
  reg [(4'ha):(1'h0)] forvar94 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg95 = (1'h0);
  reg [(5'h14):(1'h0)] reg96 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg97 = (1'h0);
  reg [(5'h10):(1'h0)] reg98 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg99 = (1'h0);
  reg [(4'hb):(1'h0)] forvar100 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg101 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg104 = (1'h0);
  reg [(4'hc):(1'h0)] reg105 = (1'h0);
  reg [(4'h8):(1'h0)] forvar106 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar110 = (1'h0);
  reg [(4'h8):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg112 = (1'h0);
  reg [(2'h3):(1'h0)] reg113 = (1'h0);
  reg [(5'h13):(1'h0)] reg114 = (1'h0);
  reg signed [(4'he):(1'h0)] reg115 = (1'h0);
  reg [(4'h8):(1'h0)] reg116 = (1'h0);
  reg [(3'h7):(1'h0)] forvar117 = (1'h0);
  reg [(5'h12):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg121 = (1'h0);
  reg [(2'h2):(1'h0)] reg122 = (1'h0);
  reg [(3'h5):(1'h0)] reg123 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg124 = (1'h0);
  reg [(5'h15):(1'h0)] forvar125 = (1'h0);
  reg [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg129 = (1'h0);
  reg [(5'h15):(1'h0)] reg130 = (1'h0);
  reg [(4'hd):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg133 = (1'h0);
  reg [(3'h6):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg135 = (1'h0);
  reg [(5'h11):(1'h0)] forvar128 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg137 = (1'h0);
  reg [(5'h15):(1'h0)] forvar138 = (1'h0);
  reg [(4'hc):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] forvar140 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg141 = (1'h0);
  reg [(2'h3):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg144 = (1'h0);
  reg [(5'h15):(1'h0)] reg145 = (1'h0);
  reg [(4'hf):(1'h0)] forvar146 = (1'h0);
  reg signed [(4'he):(1'h0)] reg147 = (1'h0);
  reg [(5'h11):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar149 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg151 = (1'h0);
  reg [(4'he):(1'h0)] reg152 = (1'h0);
  reg [(4'hc):(1'h0)] reg153 = (1'h0);
  reg [(4'h8):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg155 = (1'h0);
  reg [(4'hf):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar154 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg157 = (1'h0);
  wire [(2'h3):(1'h0)] wire158;
  wire [(3'h7):(1'h0)] wire324;
  wire signed [(4'hc):(1'h0)] wire534;
  assign y = {wire556,
                 wire555,
                 wire554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 forvar548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 forvar543,
                 reg542,
                 reg541,
                 reg540,
                 forvar539,
                 forvar538,
                 reg537,
                 reg536,
                 reg56,
                 forvar57,
                 reg58,
                 reg59,
                 reg60,
                 reg61,
                 reg62,
                 forvar63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 forvar68,
                 reg69,
                 reg70,
                 reg71,
                 reg57,
                 forvar58,
                 forvar72,
                 forvar73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 reg78,
                 reg79,
                 reg80,
                 reg81,
                 forvar82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 forvar88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 forvar93,
                 forvar94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 forvar100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 forvar106,
                 reg107,
                 reg108,
                 reg109,
                 forvar110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 forvar117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 forvar125,
                 reg126,
                 reg127,
                 reg128,
                 reg129,
                 reg130,
                 reg131,
                 forvar132,
                 reg133,
                 reg134,
                 reg135,
                 forvar128,
                 reg136,
                 reg137,
                 forvar138,
                 reg139,
                 forvar140,
                 reg141,
                 reg142,
                 reg143,
                 reg144,
                 reg145,
                 forvar146,
                 reg147,
                 reg148,
                 forvar149,
                 reg150,
                 reg151,
                 reg152,
                 reg153,
                 reg154,
                 reg155,
                 reg156,
                 forvar154,
                 reg157,
                 wire158,
                 wire324,
                 wire534,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg56 = wire53;
      if ((8'h9c))
        begin
          for (forvar57 = (1'h0); (forvar57 < (1'h1)); forvar57 = (forvar57 + (1'h1)))
            begin
              reg58 = $signed((8'ha5));
              reg59 <= (|$unsigned(reg56[(4'h8):(4'h8)]));
            end
          if (reg56)
            begin
              reg60 = "M";
              reg61 <= (^~(((~^{wire53, wire55}) ~^ reg58) ?
                  (-$signed(reg60)) : {forvar57[(1'h0):(1'h0)]}));
              reg62 <= $signed((^~wire55[(4'ha):(3'h5)]));
            end
          else
            begin
              reg60 = reg56;
              reg61 = ($signed((~&$unsigned((~&(8'ha0))))) << $signed((~|$unsigned((reg56 ?
                  forvar57 : reg61)))));
            end
          for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
            begin
              reg64 = $unsigned($signed(forvar63));
              reg65 = (({$unsigned({reg60})} ?
                      $signed(forvar63[(3'h7):(2'h2)]) : reg62) ?
                  $signed((reg59 ?
                      ((wire53 >> reg59) ?
                          (reg61 ^ reg58) : wire53[(3'h6):(2'h2)]) : (^(reg58 >>> reg60)))) : {$unsigned(($unsigned((8'haf)) + (forvar63 <<< reg61)))});
              reg66 <= $signed((((&$unsigned(reg64)) <<< $signed($signed(reg59))) || $signed($signed($unsigned(reg61)))));
              reg67 <= $unsigned(reg62[(4'hb):(1'h1)]);
            end
          for (forvar68 = (1'h0); (forvar68 < (2'h3)); forvar68 = (forvar68 + (1'h1)))
            begin
              reg69 <= (reg66[(1'h1):(1'h1)] + $unsigned(reg67));
              reg70 = (reg60 ?
                  (^~(~&((^(8'hb0)) ^ $unsigned((8'ha4))))) : (~^($unsigned("47Fgv6VvJ") ?
                      forvar68 : (forvar57 ? {reg56, forvar57} : (-wire52)))));
            end
          reg71 = forvar68;
        end
      else
        begin
          reg57 = ({$signed((forvar63 ? (^~(8'hae)) : (~&wire54))),
              forvar68[(4'h8):(1'h0)]} ^~ $unsigned(reg70));
          for (forvar58 = (1'h0); (forvar58 < (3'h4)); forvar58 = (forvar58 + (1'h1)))
            begin
              reg59 = $unsigned((wire54 == ((8'hba) ? (8'hb7) : wire53)));
              reg60 <= $unsigned(((^$signed((^~wire54))) ?
                  {$unsigned({forvar58}),
                      (~|(-reg67))} : (forvar63[(4'h8):(3'h5)] - ($unsigned(forvar57) ?
                      $signed(reg57) : $unsigned(reg60)))));
            end
          reg61 = $signed((7'h42));
          reg62 <= ($unsigned($signed($unsigned(reg66[(3'h5):(2'h3)]))) ?
              (wire54[(2'h3):(2'h3)] ?
                  {reg67[(3'h4):(1'h1)],
                      (~|(reg71 ?
                          reg65 : forvar68))} : {((7'h41) | reg69[(3'h5):(2'h3)]),
                      ((reg65 || reg58) ?
                          $unsigned(wire55) : reg65)}) : reg56[(1'h1):(1'h0)]);
        end
      for (forvar72 = (1'h0); (forvar72 < (2'h2)); forvar72 = (forvar72 + (1'h1)))
        begin
          for (forvar73 = (1'h0); (forvar73 < (1'h1)); forvar73 = (forvar73 + (1'h1)))
            begin
              reg74 <= $signed("JakZ3VzVa2bJML7bh");
              reg75 = $signed($signed((((~&forvar58) <<< $signed(reg56)) ?
                  reg62[(3'h6):(2'h2)] : (+((8'ha3) ? reg67 : wire53)))));
            end
          reg76 <= forvar58[(4'h8):(4'h8)];
          if ($unsigned(($signed(forvar73[(5'h10):(5'h10)]) ?
              {{"5qE8Z7BLmDP1", $signed(reg71)},
                  (8'ha9)} : forvar63[(2'h2):(2'h2)])))
            begin
              reg77 <= (8'hbb);
              reg78 = reg71[(3'h6):(3'h6)];
              reg79 <= forvar72;
              reg80 = reg64;
            end
          else
            begin
              reg77 = reg76[(5'h12):(5'h11)];
              reg78 = $signed($signed($signed(reg77[(2'h2):(1'h1)])));
              reg79 <= (~|reg60);
              reg80 = {forvar68[(2'h3):(1'h0)], reg76};
              reg81 = {(~^reg67)};
            end
          for (forvar82 = (1'h0); (forvar82 < (1'h1)); forvar82 = (forvar82 + (1'h1)))
            begin
              reg83 <= $signed(reg65[(2'h3):(1'h1)]);
              reg84 = reg59;
              reg85 <= $unsigned((wire53[(4'h8):(2'h3)] && (-(8'h9c))));
              reg86 = $unsigned((reg57[(4'h9):(1'h0)] ?
                  (({reg74, forvar73} <<< reg65) ?
                      reg65[(3'h5):(2'h2)] : (-(reg85 ?
                          forvar72 : reg81))) : (~&($signed(reg70) ~^ reg79))));
              reg87 = {(8'had),
                  (((~&(reg77 || reg84)) ?
                          $signed((!forvar63)) : ((~reg81) ?
                              reg83 : $unsigned(wire53))) ?
                      $unsigned(forvar68[(2'h3):(1'h1)]) : ($signed($signed(reg84)) || $unsigned((+reg62))))};
            end
          for (forvar88 = (1'h0); (forvar88 < (2'h2)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 <= ({{$signed($unsigned((8'hb3)))}} <<< forvar72[(1'h1):(1'h0)]);
              reg90 = $unsigned(((((~reg81) ^ forvar82) ?
                  reg67 : forvar88[(1'h1):(1'h0)]) > (~^(wire54[(2'h3):(1'h1)] ?
                  (reg69 ? reg76 : reg79) : $signed(reg62)))));
              reg91 <= (reg90[(4'hb):(4'h9)] ~^ ((|{"Z8xZI3ni3z",
                  reg59[(1'h0):(1'h0)]}) && $signed(($unsigned(reg65) >> (reg67 ?
                  reg83 : reg74)))));
              reg92 <= $signed(($unsigned((reg59[(2'h2):(2'h2)] ?
                  reg86 : (reg86 ?
                      (8'ha5) : reg58))) - $unsigned(forvar57[(2'h2):(1'h0)])));
            end
        end
      for (forvar93 = (1'h0); (forvar93 < (3'h4)); forvar93 = (forvar93 + (1'h1)))
        begin
          for (forvar94 = (1'h0); (forvar94 < (3'h4)); forvar94 = (forvar94 + (1'h1)))
            begin
              reg95 <= (reg76 ?
                  (~&$unsigned($unsigned((reg67 ?
                      reg58 : forvar68)))) : (($signed((&reg57)) ?
                      $signed("w") : ({reg77} - (~|reg70))) < reg77[(3'h6):(2'h2)]));
              reg96 <= $unsigned({$signed(reg58[(4'hb):(3'h6)])});
              reg97 <= ((forvar94 > ($unsigned($unsigned(reg75)) <= $signed({forvar58,
                  reg71}))) << {reg59[(3'h5):(3'h5)], {$signed((~reg62))}});
              reg98 <= (|$unsigned(reg77[(3'h4):(2'h2)]));
            end
          reg99 = ("tpKuN" ~^ $unsigned({($unsigned(reg75) > (^~reg64)),
              ("xZKhoCRSTeC2MGY" || forvar73)}));
          for (forvar100 = (1'h0); (forvar100 < (2'h2)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 <= ($unsigned(reg56[(1'h0):(1'h0)]) >= $unsigned(((8'ha9) ?
                  (^~$signed(reg67)) : ((forvar63 ? reg81 : forvar73) ?
                      reg90 : reg74[(1'h0):(1'h0)]))));
              reg102 = (~&(^~({(8'ha5), reg97} ~^ (-$signed(reg57)))));
              reg103 <= $signed(({(-$signed(forvar93))} == $unsigned($signed(((8'hbe) ?
                  reg81 : (8'hb2))))));
              reg104 <= reg87[(1'h1):(1'h0)];
              reg105 <= $unsigned((!$unsigned((reg89 ? reg97 : reg92))));
            end
          for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 <= $signed($signed({($unsigned(reg102) != ((8'hb4) * (8'h9d))),
                  $unsigned(reg96)}));
              reg108 <= reg77[(2'h3):(2'h3)];
              reg109 <= $signed((($signed(reg89) << reg97[(2'h2):(2'h2)]) ?
                  (8'hb3) : ($unsigned($signed(forvar88)) * $unsigned($unsigned(reg92)))));
            end
          for (forvar110 = (1'h0); (forvar110 < (2'h3)); forvar110 = (forvar110 + (1'h1)))
            begin
              reg111 <= reg81[(3'h7):(3'h5)];
              reg112 <= (~(|((~^(~^(8'h9c))) - $unsigned((^~reg89)))));
              reg113 <= $unsigned({forvar63[(4'hb):(2'h2)]});
              reg114 = ($unsigned(reg60) ^~ reg105);
              reg115 <= $unsigned(({$unsigned((~|reg57)),
                  (~(^~reg78))} ^~ $signed((~&"ZNkGvHJ9GBGD7"))));
            end
        end
      reg116 = (((~^$signed(reg103[(4'hd):(1'h0)])) == $signed(reg64[(3'h5):(3'h5)])) + (!($signed($signed(forvar93)) ?
          reg67 : (&(reg84 ? reg105 : reg111)))));
    end
  always
    @(posedge clk) begin
      for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
        begin
          reg118 <= reg74[(3'h5):(3'h5)];
          if ({(($unsigned((~&reg115)) ^ $signed(((8'hbc) == reg115))) || reg104[(2'h3):(1'h0)])})
            begin
              reg119 <= (reg67[(3'h5):(1'h1)] ?
                  (($signed(reg107) ?
                      forvar68[(1'h0):(1'h0)] : reg69[(4'h8):(3'h6)]) <= reg109) : {$signed($signed("wAEAN5HSqo6iyaCpP")),
                      (~$unsigned($signed(reg78)))});
              reg120 = $signed((($signed(reg83[(1'h1):(1'h1)]) < (+reg97[(2'h2):(1'h0)])) != reg59));
              reg121 = ($unsigned(((~reg91) ?
                      reg84[(2'h3):(2'h2)] : reg105[(4'h8):(3'h4)])) ?
                  reg89 : forvar57[(3'h5):(2'h2)]);
              reg122 = (($unsigned($unsigned((8'ha2))) ?
                  (~|(-reg67[(3'h7):(1'h1)])) : (~forvar68)) ^~ (&reg120));
            end
          else
            begin
              reg119 <= "aZdo3nw27";
              reg120 <= ((!((+(~^reg119)) <<< ((!reg56) | forvar82))) ^~ $unsigned((|(forvar57 == wire52[(4'he):(2'h3)]))));
              reg121 = forvar73;
              reg122 = (reg112[(3'h4):(1'h0)] - (+(~&(reg107 & reg96))));
              reg123 <= ($signed((!((reg69 > (8'ha7)) != wire54))) ?
                  ((^~((reg109 ? reg111 : reg91) >> (reg109 ?
                      reg84 : reg59))) && reg111) : ((-$signed((forvar117 ?
                      reg85 : reg87))) < reg115[(3'h6):(2'h2)]));
            end
          reg124 <= $signed((!{(~$signed(wire53)),
              (reg89 ? {reg113} : (-(8'hb2)))}));
        end
      if ($unsigned($unsigned($signed(($unsigned(reg85) ?
          reg120[(4'h9):(2'h2)] : (^reg87))))))
        begin
          for (forvar125 = (1'h0); (forvar125 < (1'h0)); forvar125 = (forvar125 + (1'h1)))
            begin
              reg126 = {(reg62[(2'h3):(1'h0)] ?
                      (8'hba) : (reg77 && (^(|reg56)))),
                  $unsigned(($unsigned((~reg114)) >>> forvar82[(1'h1):(1'h1)]))};
              reg127 = ($unsigned((reg114[(4'h9):(4'h8)] > $unsigned((forvar110 == (8'hab))))) ?
                  (reg90 ?
                      reg101[(3'h6):(2'h3)] : $signed((reg119[(4'hb):(3'h5)] ?
                          (^~reg97) : forvar82))) : $unsigned((reg95[(1'h0):(1'h0)] ?
                      $signed($unsigned(reg79)) : reg75[(2'h3):(1'h1)])));
              reg128 = forvar73[(4'hd):(4'hc)];
              reg129 = (&(~&(8'hbf)));
            end
          reg130 <= (&reg56);
          reg131 = (forvar73 ^~ reg56);
          for (forvar132 = (1'h0); (forvar132 < (1'h0)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= (($signed(($unsigned(reg69) ?
                          $unsigned(reg89) : reg76)) ?
                      $signed($unsigned((forvar110 ~^ reg97))) : reg123) ?
                  $signed(reg84) : reg118[(4'h9):(3'h7)]);
              reg134 <= $signed(forvar117[(3'h4):(1'h1)]);
            end
          if ($unsigned(((^wire54) & reg80)))
            begin
              reg135 = (!{((((8'haa) < (8'ha7)) >= (reg119 ?
                      reg89 : wire55)) || ($signed(reg118) ?
                      (~forvar106) : (reg60 != (8'h9d)))),
                  reg105[(3'h5):(3'h4)]});
            end
          else
            begin
              reg135 = {$unsigned($unsigned(forvar58))};
            end
        end
      else
        begin
          for (forvar125 = (1'h0); (forvar125 < (2'h3)); forvar125 = (forvar125 + (1'h1)))
            begin
              reg126 <= reg69[(4'h8):(3'h6)];
              reg127 <= ((|(({reg119} || (~&reg91)) ?
                  reg103 : ((reg64 == reg127) != $unsigned(reg127)))) != (((8'hbc) ?
                      ((-reg95) ? reg99 : reg134) : {$unsigned(reg131)}) ?
                  reg58[(4'h9):(3'h4)] : $signed(((forvar72 <= (8'hb6)) | forvar100[(3'h5):(1'h1)]))));
            end
          for (forvar128 = (1'h0); (forvar128 < (1'h1)); forvar128 = (forvar128 + (1'h1)))
            begin
              reg129 <= reg76;
              reg130 = $signed((8'haf));
              reg131 <= {$unsigned($signed(forvar63[(2'h3):(1'h0)]))};
            end
        end
      reg136 <= $unsigned($signed($unsigned(wire52[(4'he):(4'h8)])));
      reg137 = reg107[(4'ha):(1'h1)];
      for (forvar138 = (1'h0); (forvar138 < (1'h1)); forvar138 = (forvar138 + (1'h1)))
        begin
          reg139 = {(reg85 ?
                  $signed(((+reg91) ?
                      (!forvar110) : (reg96 != reg112))) : $signed($signed(reg130))),
              $signed(((+$unsigned(reg113)) ?
                  (~|(reg120 ? reg64 : forvar82)) : $unsigned((~|reg95))))};
          for (forvar140 = (1'h0); (forvar140 < (1'h1)); forvar140 = (forvar140 + (1'h1)))
            begin
              reg141 <= (($signed((&"0YRVXOdlB")) * reg69) ?
                  $signed(((reg107 > (7'h43)) >> $unsigned({reg109,
                      reg69}))) : (^~reg58[(4'hc):(4'hb)]));
            end
          if (forvar68[(4'hc):(3'h7)])
            begin
              reg142 <= $signed($unsigned($unsigned((&$signed(forvar100)))));
              reg143 = (forvar128[(1'h0):(1'h0)] ?
                  $unsigned(reg67[(3'h4):(1'h1)]) : $unsigned((~&(+(8'hae)))));
            end
          else
            begin
              reg142 <= ((+$signed($unsigned($unsigned(reg120)))) ^ forvar93[(4'he):(3'h4)]);
              reg143 = $unsigned(reg66);
              reg144 = ((reg78[(5'h10):(4'hd)] > "86npJbqn9OqkDqkh") & forvar132[(4'h9):(2'h3)]);
              reg145 <= $unsigned($unsigned(($unsigned(wire52[(4'hc):(2'h3)]) ?
                  ($unsigned(reg92) | {reg126}) : (~reg109[(2'h2):(1'h1)]))));
            end
          for (forvar146 = (1'h0); (forvar146 < (2'h2)); forvar146 = (forvar146 + (1'h1)))
            begin
              reg147 = forvar138[(4'h8):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ((~^((((forvar72 & reg104) - reg119[(5'h14):(2'h3)]) > ($unsigned(reg133) ~^ (7'h44))) * $signed(({reg81,
              reg126} ?
          $unsigned(reg133) : reg124)))))
        begin
          reg148 <= $signed(({{(8'ha5)}} ^ reg121[(1'h1):(1'h1)]));
          for (forvar149 = (1'h0); (forvar149 < (1'h1)); forvar149 = (forvar149 + (1'h1)))
            begin
              reg150 <= ((8'hbc) ?
                  reg98 : $signed((reg144[(4'hb):(1'h1)] ?
                      (!(forvar58 != reg147)) : $unsigned((forvar63 * (8'hb8))))));
              reg151 = (reg139 ?
                  ("LqN" < $signed(((reg143 ?
                      reg61 : (8'h9d)) >= $signed(reg86)))) : $signed(reg143));
              reg152 <= (~&((+(forvar73 << (forvar128 ^ reg112))) ?
                  {$signed(((8'hb6) != reg70)),
                      ((7'h43) ?
                          (|reg145) : reg123[(3'h4):(2'h2)])} : $unsigned((~(reg81 ?
                      reg119 : (8'ha7))))));
              reg153 = ((+{(|(reg120 ?
                      (7'h41) : reg64))}) <= $signed(($signed(reg136[(2'h2):(1'h1)]) ?
                  $unsigned(((8'hba) <= reg59)) : (-reg126[(3'h4):(2'h3)]))));
            end
          if ($unsigned($unsigned((~&reg97))))
            begin
              reg154 <= $signed($unsigned(("aJlABHE" ?
                  $signed($unsigned(reg134)) : reg131)));
            end
          else
            begin
              reg154 = (&$unsigned($unsigned(reg76)));
            end
          reg155 <= ($unsigned($signed((reg104 ?
              {reg144} : (reg127 && reg90)))) || (~|(-reg123[(3'h5):(1'h0)])));
          reg156 = reg115;
        end
      else
        begin
          reg148 <= "OsDol6MXKkd";
          for (forvar149 = (1'h0); (forvar149 < (1'h0)); forvar149 = (forvar149 + (1'h1)))
            begin
              reg150 = ($unsigned($signed({$unsigned(reg129),
                      $signed(reg56)})) ?
                  reg85 : ({((+reg78) > (reg112 ? wire54 : reg145)),
                          $signed(reg108)} ?
                      {reg89} : ({$unsigned(reg147)} >>> ($signed((8'haf)) | $signed(reg143)))));
              reg151 <= $unsigned((8'hb8));
              reg152 = reg156;
              reg153 <= (~(7'h40));
            end
          for (forvar154 = (1'h0); (forvar154 < (2'h2)); forvar154 = (forvar154 + (1'h1)))
            begin
              reg155 = ((reg87 ?
                  forvar72 : (((reg152 ? reg130 : forvar68) ^~ (8'hb8)) ?
                      reg145[(3'h5):(3'h5)] : "EUk6qRe9kW")) * (!(!($signed(reg91) ?
                  (reg67 ? reg151 : reg150) : $signed(reg153)))));
              reg156 <= reg104;
              reg157 <= (~^reg120[(5'h12):(3'h6)]);
            end
        end
    end
  assign wire158 = $unsigned((|(|{((8'ha7) ? (8'hb7) : forvar93)})));
  module159 modinst325 (.wire162(reg74), .clk(clk), .wire161(reg67), .wire160(forvar128), .wire163(forvar57), .y(wire324));
  module326 modinst535 (.wire328(reg156), .clk(clk), .wire327(forvar146), .wire329(reg133), .wire330(reg152), .y(wire534), .wire331(reg57));
  always
    @(posedge clk) begin
      reg536 = $signed((wire52[(4'he):(4'ha)] ? reg145 : reg76[(4'hb):(4'hb)]));
      reg537 <= $unsigned(($signed((~|$signed(reg78))) >> (($signed(reg80) && reg152) ?
          ((8'hac) ^ (reg97 * reg103)) : $unsigned($unsigned(reg86)))));
      for (forvar538 = (1'h0); (forvar538 < (1'h0)); forvar538 = (forvar538 + (1'h1)))
        begin
          for (forvar539 = (1'h0); (forvar539 < (3'h4)); forvar539 = (forvar539 + (1'h1)))
            begin
              reg540 <= reg155[(2'h2):(2'h2)];
              reg541 = (((~^reg144) >> ($signed(reg78) ?
                      (8'hb5) : ($unsigned(reg79) ? $signed(reg70) : reg147))) ?
                  $signed((&$signed(reg59[(2'h3):(2'h2)]))) : ("L4mRSKYzxsgpATzOUo" ~^ ((reg154 ?
                          (reg107 ? (8'ha9) : (7'h42)) : reg92[(3'h6):(1'h1)]) ?
                      {{reg113}} : reg121[(4'h8):(3'h5)])));
              reg542 = $signed($signed(($unsigned((forvar73 ?
                      forvar132 : reg95)) ?
                  reg131 : (|$signed((8'hb3))))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg87)
        begin
          for (forvar543 = (1'h0); (forvar543 < (1'h0)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 = $signed("Dtsx7AVzd92Rfxg");
              reg545 <= $unsigned(reg145[(2'h2):(2'h2)]);
              reg546 = forvar138;
            end
        end
      else
        begin
          for (forvar543 = (1'h0); (forvar543 < (1'h0)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 = reg145;
              reg545 = (~^((reg136 != (8'hbe)) ? wire52 : reg131));
              reg546 <= reg89;
              reg547 = (((reg143[(3'h4):(1'h0)] & (reg116[(2'h2):(2'h2)] ?
                          (reg103 >>> (8'h9e)) : "zBsUfd7C6ra")) ?
                      (reg77 >= $signed((reg118 ?
                          reg111 : reg111))) : forvar140[(1'h1):(1'h1)]) ?
                  reg145[(1'h0):(1'h0)] : (8'haa));
            end
          for (forvar548 = (1'h0); (forvar548 < (3'h4)); forvar548 = (forvar548 + (1'h1)))
            begin
              reg549 = $unsigned($signed((8'hb0)));
              reg550 = reg114[(2'h3):(2'h2)];
            end
          reg551 <= reg128[(4'h9):(4'h8)];
          reg552 <= $unsigned((($unsigned((~^reg103)) ?
              ((reg542 << reg151) ?
                  {reg541,
                      (8'hb1)} : $signed(wire52)) : {reg77}) == (~^$unsigned({forvar140,
              reg134}))));
        end
      reg553 = ($signed($unsigned(reg549[(2'h3):(2'h2)])) ?
          (~&reg57) : $signed(reg143));
    end
  assign wire554 = (^$unsigned(wire53[(5'h11):(5'h11)]));
  assign wire555 = {reg550[(4'hd):(1'h1)], $unsigned(reg60)};
  assign wire556 = (forvar539 ?
                       ((($unsigned(forvar73) <<< (reg56 ?
                               wire54 : (8'hae))) & reg111) ?
                           $signed($signed((forvar93 * reg153))) : (-({(8'hb6),
                               forvar128} - reg540[(3'h5):(3'h5)]))) : (^~$signed((reg78[(2'h2):(2'h2)] == ((7'h40) ^~ reg84)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module326
#( parameter param532 = (((~(((8'ha5) >> (8'hb1)) ? ((8'ha0) ? (8'ha1) : (8'h9f)) : ((8'hbc) ? (8'hb0) : (8'hb1)))) ^~ ((~{(8'hb4)}) < ({(8'ha1)} >= ((8'ha7) >>> (8'ha5))))) - ((~^(8'h9d)) ? ((&(7'h42)) + ((-(8'h9c)) ? ((8'haf) ? (8'h9d) : (8'ha8)) : ((8'hb4) <<< (8'haf)))) : (((~|(8'ha8)) ? (~&(8'hb6)) : (^(8'hab))) << (~|(~|(8'ha7))))))
, parameter param533 = param532 )
(y, clk, wire331, wire330, wire329, wire328, wire327);
  output wire [(32'h899):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire331;
  input wire [(4'h8):(1'h0)] wire330;
  input wire [(4'ha):(1'h0)] wire329;
  input wire signed [(4'hf):(1'h0)] wire328;
  input wire signed [(4'ha):(1'h0)] wire327;
  wire [(4'h8):(1'h0)] wire531;
  wire [(5'h11):(1'h0)] wire530;
  reg signed [(5'h11):(1'h0)] reg529 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar528 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg526 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg524 = (1'h0);
  reg [(4'hf):(1'h0)] forvar521 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg523 = (1'h0);
  reg [(5'h12):(1'h0)] reg522 = (1'h0);
  reg [(4'hf):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar520 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg519 = (1'h0);
  reg [(3'h4):(1'h0)] reg518 = (1'h0);
  reg [(2'h3):(1'h0)] reg517 = (1'h0);
  reg [(3'h7):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg515 = (1'h0);
  reg [(3'h4):(1'h0)] forvar514 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg511 = (1'h0);
  reg [(5'h12):(1'h0)] reg510 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg509 = (1'h0);
  reg [(4'hd):(1'h0)] reg508 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg506 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg504 = (1'h0);
  reg [(4'he):(1'h0)] reg503 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar501 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg499 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg498 = (1'h0);
  reg [(4'hd):(1'h0)] reg497 = (1'h0);
  reg [(4'ha):(1'h0)] reg496 = (1'h0);
  reg [(5'h15):(1'h0)] forvar495 = (1'h0);
  reg [(5'h15):(1'h0)] reg494 = (1'h0);
  reg [(5'h10):(1'h0)] reg493 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar492 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg491 = (1'h0);
  reg [(4'hd):(1'h0)] forvar490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg489 = (1'h0);
  reg [(3'h5):(1'h0)] forvar488 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg487 = (1'h0);
  reg [(5'h10):(1'h0)] reg486 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg484 = (1'h0);
  reg signed [(4'he):(1'h0)] reg483 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg [(5'h12):(1'h0)] forvar480 = (1'h0);
  reg [(5'h14):(1'h0)] reg479 = (1'h0);
  reg [(3'h5):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar474 = (1'h0);
  wire [(3'h4):(1'h0)] wire473;
  reg signed [(4'hc):(1'h0)] reg472 = (1'h0);
  reg [(4'hc):(1'h0)] reg471 = (1'h0);
  reg [(3'h6):(1'h0)] reg470 = (1'h0);
  reg [(4'hd):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg468 = (1'h0);
  reg [(3'h7):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar466 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar465 = (1'h0);
  reg [(2'h3):(1'h0)] reg464 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg463 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg462 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg461 = (1'h0);
  reg [(5'h14):(1'h0)] reg460 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar459 = (1'h0);
  reg [(5'h13):(1'h0)] reg458 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg457 = (1'h0);
  reg [(5'h10):(1'h0)] reg456 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg455 = (1'h0);
  reg [(2'h2):(1'h0)] reg454 = (1'h0);
  reg [(5'h11):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar451 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg450 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg449 = (1'h0);
  reg [(4'he):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar447 = (1'h0);
  reg [(3'h5):(1'h0)] forvar446 = (1'h0);
  wire [(4'h8):(1'h0)] wire445;
  reg [(4'ha):(1'h0)] reg444 = (1'h0);
  reg [(4'he):(1'h0)] reg443 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg442 = (1'h0);
  reg [(4'ha):(1'h0)] reg441 = (1'h0);
  reg [(3'h5):(1'h0)] reg440 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg439 = (1'h0);
  reg [(3'h4):(1'h0)] reg438 = (1'h0);
  reg [(3'h5):(1'h0)] reg437 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg436 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg435 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg433 = (1'h0);
  reg [(4'hb):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg431 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar430 = (1'h0);
  reg [(5'h14):(1'h0)] reg429 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg428 = (1'h0);
  reg [(5'h10):(1'h0)] reg427 = (1'h0);
  reg [(5'h12):(1'h0)] forvar426 = (1'h0);
  reg [(5'h15):(1'h0)] reg425 = (1'h0);
  reg [(2'h2):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg422 = (1'h0);
  reg [(4'ha):(1'h0)] forvar421 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg420 = (1'h0);
  reg [(4'hd):(1'h0)] reg419 = (1'h0);
  reg [(4'h8):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar417 = (1'h0);
  reg [(3'h4):(1'h0)] reg416 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar415 = (1'h0);
  reg [(5'h12):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg410 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg408 = (1'h0);
  reg [(4'h8):(1'h0)] reg407 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg406 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg405 = (1'h0);
  reg [(3'h6):(1'h0)] forvar404 = (1'h0);
  reg [(5'h14):(1'h0)] forvar403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg402 = (1'h0);
  wire [(4'hb):(1'h0)] wire401;
  reg [(5'h15):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg399 = (1'h0);
  reg [(4'hf):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg397 = (1'h0);
  reg [(5'h12):(1'h0)] forvar396 = (1'h0);
  reg [(5'h11):(1'h0)] reg395 = (1'h0);
  reg [(4'hd):(1'h0)] reg394 = (1'h0);
  reg [(3'h7):(1'h0)] reg393 = (1'h0);
  reg [(5'h15):(1'h0)] reg392 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg391 = (1'h0);
  reg [(5'h15):(1'h0)] forvar390 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar389 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg388 = (1'h0);
  reg [(5'h14):(1'h0)] reg387 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg385 = (1'h0);
  reg [(4'ha):(1'h0)] reg384 = (1'h0);
  reg [(5'h13):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg382 = (1'h0);
  reg [(2'h3):(1'h0)] reg381 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar377 = (1'h0);
  reg [(2'h2):(1'h0)] reg376 = (1'h0);
  reg [(2'h2):(1'h0)] reg375 = (1'h0);
  reg [(4'hc):(1'h0)] reg374 = (1'h0);
  reg [(4'hd):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar372 = (1'h0);
  reg [(4'h8):(1'h0)] reg371 = (1'h0);
  reg [(3'h4):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg368 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg367 = (1'h0);
  reg [(4'h8):(1'h0)] reg366 = (1'h0);
  reg [(2'h2):(1'h0)] forvar365 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar364 = (1'h0);
  reg [(5'h12):(1'h0)] reg363 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg362 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg361 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar360 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg359 = (1'h0);
  reg [(5'h10):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar357 = (1'h0);
  reg [(2'h3):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg355 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar354 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar353 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg352 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg351 = (1'h0);
  wire [(4'h8):(1'h0)] wire350;
  wire signed [(4'h8):(1'h0)] wire349;
  reg [(5'h10):(1'h0)] reg348 = (1'h0);
  reg [(2'h3):(1'h0)] reg347 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar346 = (1'h0);
  reg [(2'h3):(1'h0)] reg345 = (1'h0);
  reg [(4'ha):(1'h0)] forvar344 = (1'h0);
  reg [(3'h7):(1'h0)] reg343 = (1'h0);
  reg [(5'h13):(1'h0)] reg342 = (1'h0);
  reg [(2'h2):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar340 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg339 = (1'h0);
  reg [(2'h2):(1'h0)] reg338 = (1'h0);
  reg [(3'h6):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar335 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire334;
  wire signed [(4'hb):(1'h0)] wire333;
  wire [(5'h11):(1'h0)] wire332;
  assign y = {wire531,
                 wire530,
                 reg529,
                 forvar528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 forvar521,
                 reg520,
                 reg523,
                 reg522,
                 reg521,
                 forvar520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 forvar495,
                 reg494,
                 reg493,
                 forvar492,
                 reg491,
                 forvar490,
                 reg489,
                 forvar488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 forvar474,
                 wire473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 forvar466,
                 forvar465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 forvar459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 forvar451,
                 reg450,
                 reg449,
                 reg448,
                 forvar447,
                 forvar446,
                 wire445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 forvar434,
                 reg433,
                 reg432,
                 reg431,
                 forvar430,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 forvar417,
                 reg416,
                 forvar415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 forvar403,
                 reg402,
                 wire401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 forvar396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 forvar390,
                 forvar389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 forvar372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 forvar365,
                 forvar364,
                 reg363,
                 reg362,
                 reg361,
                 forvar360,
                 reg359,
                 reg358,
                 forvar357,
                 reg356,
                 reg355,
                 forvar354,
                 forvar353,
                 reg352,
                 reg351,
                 wire350,
                 wire349,
                 reg348,
                 reg347,
                 forvar346,
                 reg345,
                 forvar344,
                 reg343,
                 reg342,
                 reg341,
                 forvar340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 forvar335,
                 wire334,
                 wire333,
                 wire332,
                 (1'h0)};
  assign wire332 = (!($signed($signed((wire330 ~^ wire327))) >> $unsigned(wire328[(1'h0):(1'h0)])));
  assign wire333 = wire327;
  assign wire334 = {$unsigned($unsigned($unsigned((!wire331))))};
  always
    @(posedge clk) begin
      for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
        begin
          if ((|($unsigned(({wire331} ?
              wire328 : $signed(wire334))) || ($unsigned("w") ?
              $signed((wire331 ?
                  forvar335 : wire330)) : $unsigned(forvar335)))))
            begin
              reg336 <= (^({$unsigned("b"),
                  wire331[(3'h6):(3'h5)]} >> (^~forvar335)));
              reg337 <= (~^($signed($signed(wire329)) < $signed(($signed(wire328) <<< $signed(wire332)))));
              reg338 <= {(~^$unsigned($unsigned((+wire332))))};
              reg339 = wire331;
            end
          else
            begin
              reg336 = $unsigned((8'ha6));
              reg337 = wire327;
              reg338 <= $unsigned({forvar335[(3'h4):(1'h1)]});
              reg339 = ("2LzeTE2SH3qIh" ?
                  (reg339 ?
                      ("Mhbs39ay7S8LXNbY" * reg338[(1'h0):(1'h0)]) : $signed((~&(^wire334)))) : $unsigned(wire332[(3'h7):(3'h5)]));
            end
          for (forvar340 = (1'h0); (forvar340 < (1'h0)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= $signed(reg336);
              reg342 = $unsigned($unsigned({($signed(reg337) ?
                      $signed(reg338) : (wire332 ? reg338 : reg337))}));
              reg343 = reg339;
            end
          for (forvar344 = (1'h0); (forvar344 < (2'h2)); forvar344 = (forvar344 + (1'h1)))
            begin
              reg345 <= "fMRGbFFV1ldYDS";
            end
          for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 <= (reg337 <<< (wire332 ?
                  (&$unsigned((^~(8'hba)))) : wire330));
              reg348 <= ($unsigned({{{wire329},
                          (reg345 ? forvar346 : reg342)}}) ?
                  (&reg336) : reg337[(1'h1):(1'h0)]);
            end
        end
    end
  assign wire349 = wire330;
  assign wire350 = (wire334 ?
                       ("JOocWAlfMiK" || (((!(8'ha7)) << reg348[(3'h7):(2'h2)]) <<< ((~|wire328) ?
                           $unsigned(reg341) : (reg339 >>> (8'hb8))))) : ($unsigned($signed(forvar346)) ?
                           (~^wire333[(2'h2):(2'h2)]) : wire334));
  always
    @(posedge clk) begin
      reg351 = (((-$signed($signed((8'ha5)))) ? (8'hbc) : wire349) ?
          (8'haa) : "QUl");
      reg352 = {$unsigned($unsigned(wire327[(4'h8):(3'h7)])),
          {wire331[(3'h4):(3'h4)],
              {((-wire329) ? $signed(reg345) : (wire329 >= reg337)),
                  {wire330, (reg337 ? reg348 : wire350)}}}};
    end
  always
    @(posedge clk) begin
      for (forvar353 = (1'h0); (forvar353 < (3'h4)); forvar353 = (forvar353 + (1'h1)))
        begin
          for (forvar354 = (1'h0); (forvar354 < (1'h0)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 <= $unsigned({$signed({"hAL88L2iiKDm0"})});
              reg356 = ({wire334,
                      ((((8'hb9) | reg351) ? {reg343} : $unsigned(reg355)) ?
                          wire331 : (7'h40))} ?
                  $unsigned(((reg341 ?
                      forvar335[(3'h4):(2'h3)] : $signed((7'h44))) < reg338[(1'h1):(1'h1)])) : reg345[(1'h0):(1'h0)]);
            end
          for (forvar357 = (1'h0); (forvar357 < (1'h0)); forvar357 = (forvar357 + (1'h1)))
            begin
              reg358 <= reg339[(3'h6):(1'h1)];
              reg359 = {$unsigned(($unsigned((~&forvar353)) ?
                      $signed(reg338) : $signed($signed(wire329))))};
            end
        end
      for (forvar360 = (1'h0); (forvar360 < (3'h4)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 = ($signed(reg347) ?
              $unsigned((-(^{wire331}))) : {reg339[(4'hd):(3'h7)],
                  $signed(reg358)});
          reg362 <= (((~&wire329[(4'h9):(1'h0)]) * $unsigned($signed(forvar360[(1'h0):(1'h0)]))) != (($signed(((7'h44) ?
                      wire331 : reg341)) ?
                  (8'ha9) : $signed($signed(forvar346))) ?
              $unsigned({(reg343 && reg342),
                  {reg348}}) : ($signed($unsigned(forvar360)) ~^ "Ji")));
          reg363 = "yHyBp1";
        end
      for (forvar364 = (1'h0); (forvar364 < (1'h1)); forvar364 = (forvar364 + (1'h1)))
        begin
          for (forvar365 = (1'h0); (forvar365 < (3'h4)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 <= forvar364[(3'h5):(1'h0)];
              reg367 = {$unsigned(forvar354[(4'h9):(3'h4)]),
                  $signed(forvar353[(2'h3):(1'h1)])};
              reg368 <= $signed(((forvar357[(3'h5):(3'h5)] >>> ({wire327,
                      forvar360} ^~ (reg338 ? wire328 : reg363))) ?
                  forvar354[(3'h7):(1'h0)] : $unsigned(((forvar353 & forvar344) <<< forvar354))));
            end
          if (({(wire332[(4'hd):(3'h4)] >>> $unsigned(reg368[(2'h2):(1'h1)]))} ?
              (wire334[(2'h2):(1'h0)] < (8'hbe)) : (7'h42)))
            begin
              reg369 <= {{{(+wire331)},
                      $signed((wire331[(1'h0):(1'h0)] ?
                          wire349 : $signed(reg368)))}};
              reg370 <= (wire330 ?
                  $signed($unsigned($signed($signed(reg351)))) : {$signed($unsigned(reg337[(3'h4):(1'h0)])),
                      wire349[(3'h4):(1'h0)]});
            end
          else
            begin
              reg369 <= $signed($unsigned(((|$unsigned((7'h42))) ?
                  ($signed(reg356) * (reg348 ?
                      reg352 : forvar354)) : $signed((+reg362)))));
              reg370 <= {((-(~(reg361 ^~ reg341))) ?
                      $unsigned(wire328) : $signed((+(reg336 ?
                          wire331 : forvar360)))),
                  reg351[(2'h2):(2'h2)]};
              reg371 = (wire328 > wire330);
            end
          for (forvar372 = (1'h0); (forvar372 < (1'h0)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 = reg356[(2'h2):(1'h0)];
              reg374 <= (((8'ha7) <= {({wire329, reg363} ?
                          (^forvar372) : (wire327 ? wire331 : forvar346)),
                      (reg342 & (8'hb9))}) ?
                  reg363 : wire350);
              reg375 = (-(-(8'hbf)));
              reg376 = reg347[(1'h0):(1'h0)];
            end
          for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 <= (|"7G");
              reg379 <= ($signed(($signed((wire328 ?
                  reg359 : (8'ha0))) ~^ $signed({(8'ha7),
                  reg368}))) << ($unsigned($unsigned((~^forvar346))) > ((reg356 ?
                  wire327[(1'h0):(1'h0)] : $signed(reg355)) << (forvar340[(4'hd):(3'h6)] ?
                  reg348 : wire349))));
              reg380 <= wire329;
            end
          reg381 = reg359;
        end
      if ((-(+wire327[(2'h2):(2'h2)])))
        begin
          if ($signed(forvar357))
            begin
              reg382 <= ((($unsigned(reg342) >>> $unsigned($unsigned(reg355))) >= $unsigned($signed(reg359))) & reg371[(3'h5):(1'h0)]);
            end
          else
            begin
              reg382 = $signed($unsigned((!$unsigned($unsigned(reg339)))));
              reg383 = $signed(((&$unsigned($unsigned(reg373))) ?
                  (!{(reg352 ? reg362 : (8'h9f)),
                      reg376}) : (reg373[(4'hc):(3'h4)] * reg373)));
              reg384 <= ($unsigned({$unsigned($signed(reg359)),
                  reg342}) <= $unsigned((8'ha3)));
              reg385 = $signed((($signed($unsigned(wire350)) * $signed($signed(reg369))) * (reg352 * {(7'h41),
                  wire334})));
            end
        end
      else
        begin
          if (forvar354)
            begin
              reg382 = $signed((+(~|{(reg352 ? reg342 : reg382), reg385})));
              reg383 = (($unsigned((|(reg345 ?
                      wire349 : wire350))) + (~&reg361[(2'h3):(1'h0)])) ?
                  ($unsigned(reg362[(1'h0):(1'h0)]) + reg384[(2'h2):(1'h1)]) : wire333[(4'h8):(3'h6)]);
              reg384 = reg382;
              reg385 = (((~(-(reg339 != reg380))) || $signed((&(^~forvar360)))) == $signed(reg366));
              reg386 = (-(-(|(+((8'hae) || reg379)))));
            end
          else
            begin
              reg382 <= (-(8'hac));
            end
          reg387 <= reg343[(1'h0):(1'h0)];
          reg388 <= $signed($signed(forvar364));
        end
      for (forvar389 = (1'h0); (forvar389 < (1'h1)); forvar389 = (forvar389 + (1'h1)))
        begin
          for (forvar390 = (1'h0); (forvar390 < (2'h3)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 = reg367[(4'hf):(2'h2)];
              reg392 <= reg378[(3'h5):(2'h3)];
              reg393 <= (-$signed((((reg370 - wire333) == (+reg387)) ?
                  $unsigned(reg358) : reg385)));
              reg394 = ((!reg362[(2'h2):(2'h2)]) > (reg393[(3'h7):(1'h0)] >= (((forvar340 >>> reg393) && $unsigned(reg359)) ?
                  {(reg358 ? forvar390 : reg339),
                      ((8'had) ? reg384 : reg381)} : reg358)));
              reg395 <= (reg381[(2'h3):(2'h2)] ~^ ((reg342 ^ $unsigned((wire333 ?
                      reg342 : wire332))) ?
                  {({(8'h9f),
                          forvar335} << "kDKTuUR7AWtnL")} : $signed((^{(8'hbf)}))));
            end
          for (forvar396 = (1'h0); (forvar396 < (3'h4)); forvar396 = (forvar396 + (1'h1)))
            begin
              reg397 = (^~$signed(forvar372));
              reg398 <= reg379[(1'h0):(1'h0)];
              reg399 <= $unsigned($unsigned({(wire329[(4'h9):(3'h7)] && "Ci7qSCG")}));
              reg400 <= reg339;
            end
        end
    end
  assign wire401 = ((!(|((7'h41) ?
                       reg358[(1'h0):(1'h0)] : $signed(reg348)))) + reg386[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg402 = forvar357;
      for (forvar403 = (1'h0); (forvar403 < (1'h0)); forvar403 = (forvar403 + (1'h1)))
        begin
          for (forvar404 = (1'h0); (forvar404 < (2'h3)); forvar404 = (forvar404 + (1'h1)))
            begin
              reg405 = $signed($unsigned((-reg392)));
              reg406 = reg348[(3'h7):(2'h3)];
              reg407 <= ($signed((~|(forvar377[(1'h1):(1'h0)] >> reg382[(4'hd):(4'h8)]))) ?
                  $signed(reg345) : $signed(($unsigned(forvar404) > ((reg359 <= wire331) ?
                      (~|reg352) : {(8'haf), wire350}))));
              reg408 <= ((+$signed({$signed(reg384)})) ? (^{reg392}) : reg339);
            end
          if ({wire331[(3'h7):(2'h2)],
              {reg341,
                  (+{(reg373 ? forvar344 : forvar403),
                      (reg337 || forvar360)})}})
            begin
              reg409 = $signed((+(($signed(wire328) ^ (forvar390 != reg392)) << ($signed(reg380) ?
                  reg392 : (^~reg369)))));
              reg410 = wire350;
              reg411 = forvar377[(2'h2):(1'h1)];
              reg412 = $signed(reg398[(2'h3):(2'h2)]);
              reg413 <= (forvar364 ?
                  (&reg337[(1'h0):(1'h0)]) : $signed($signed(forvar346[(2'h2):(1'h0)])));
            end
          else
            begin
              reg409 = $unsigned($signed(reg394));
              reg410 = wire334[(1'h0):(1'h0)];
              reg411 <= ((($signed(wire349[(2'h2):(1'h1)]) >> reg410[(4'h8):(3'h5)]) ~^ (-reg359)) && (-reg402[(4'h8):(3'h7)]));
              reg412 <= (~forvar346[(2'h2):(1'h0)]);
            end
          reg414 <= (($unsigned((|(reg369 ? reg359 : forvar344))) ?
              {wire349,
                  (|$unsigned(reg361))} : (^~("pZ" * wire328))) ~^ (!($unsigned($unsigned(wire349)) ?
              ($signed((8'h9d)) ?
                  reg336[(3'h4):(2'h3)] : (reg376 && reg366)) : {(wire349 ~^ reg381),
                  $unsigned(wire349)})));
          for (forvar415 = (1'h0); (forvar415 < (1'h0)); forvar415 = (forvar415 + (1'h1)))
            begin
              reg416 = $unsigned($signed($unsigned(reg352[(2'h2):(1'h1)])));
            end
          for (forvar417 = (1'h0); (forvar417 < (3'h4)); forvar417 = (forvar417 + (1'h1)))
            begin
              reg418 <= ((-(-$signed((&reg352)))) << (reg373 - wire327[(4'h9):(3'h6)]));
              reg419 = (&(($signed($unsigned((8'h9c))) | $unsigned((reg371 ?
                      reg409 : reg397))) ?
                  $signed(({reg394} ?
                      forvar404 : (reg347 ?
                          reg355 : (8'hbf)))) : reg402[(1'h0):(1'h0)]));
              reg420 <= (8'ha5);
            end
        end
      for (forvar421 = (1'h0); (forvar421 < (2'h2)); forvar421 = (forvar421 + (1'h1)))
        begin
          if (($unsigned({($signed((8'hb0)) ?
                  $unsigned(reg384) : $unsigned(reg384))}) <<< (($signed((~forvar340)) ?
                  {reg392} : (~&(forvar417 != (8'hb1)))) ?
              (~|(~{(8'h9d)})) : {((^~reg384) ? (-reg368) : $signed(wire349)),
                  reg398})))
            begin
              reg422 <= $signed("g1zNDfEFFPZzh7mhtqTp");
              reg423 = (reg402[(3'h4):(1'h1)] << (((8'hab) ?
                  ((&reg339) ?
                      (^~reg375) : reg343) : reg338[(2'h2):(2'h2)]) >>> (($unsigned(wire327) ?
                  $unsigned(forvar389) : $unsigned((8'hac))) ^ $unsigned({(8'hae)}))));
              reg424 <= (reg385 == ($unsigned(reg356[(1'h1):(1'h0)]) != ((reg405 ?
                      $unsigned(reg339) : {reg409}) ?
                  $unsigned((reg386 != wire332)) : (|{wire401, reg393}))));
              reg425 = (!$signed(reg413));
            end
          else
            begin
              reg422 <= ($unsigned($unsigned(($unsigned(reg345) ?
                  $unsigned(reg374) : reg399))) >= (|(((reg424 ?
                          reg375 : (8'hb1)) ?
                      (~|reg368) : forvar417[(4'h9):(4'h9)]) ?
                  reg384[(2'h3):(1'h0)] : $unsigned((|reg402)))));
              reg423 <= {((~^reg370[(3'h4):(1'h0)]) != $signed((|(|reg410))))};
              reg424 = reg418[(3'h5):(1'h1)];
            end
          for (forvar426 = (1'h0); (forvar426 < (2'h3)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 <= $signed((~|((^~(reg388 ? forvar389 : wire349)) ?
                  $signed($unsigned(forvar417)) : $unsigned((8'hab)))));
              reg428 = $unsigned((-forvar403[(5'h13):(5'h10)]));
              reg429 <= {$signed(($signed((^~wire328)) & ((^~(8'ha6)) ?
                      forvar364 : (+forvar344)))),
                  $signed(((((8'hb2) ?
                          reg361 : forvar353) ^ (forvar360 >= reg412)) ?
                      $signed($signed((8'ha1))) : (+$unsigned(reg352))))};
            end
          for (forvar430 = (1'h0); (forvar430 < (1'h0)); forvar430 = (forvar430 + (1'h1)))
            begin
              reg431 = reg367[(1'h1):(1'h1)];
              reg432 <= {(8'hb5)};
            end
        end
      reg433 = $signed($signed({(reg362[(2'h3):(1'h0)] ?
              forvar344[(2'h2):(2'h2)] : ((8'ha5) <= reg399))}));
      for (forvar434 = (1'h0); (forvar434 < (2'h2)); forvar434 = (forvar434 + (1'h1)))
        begin
          reg435 <= reg342[(1'h1):(1'h1)];
          if ($signed(($signed(reg406[(1'h1):(1'h0)]) ?
              $unsigned($signed((~&reg388))) : $signed($unsigned($signed(reg337))))))
            begin
              reg436 <= $signed((+forvar340[(4'hc):(2'h2)]));
              reg437 <= ({reg339[(4'hf):(2'h3)],
                  reg402[(3'h6):(2'h2)]} <= (~|$signed($signed(forvar421[(4'ha):(4'h9)]))));
            end
          else
            begin
              reg436 <= reg385;
              reg437 = (!{(forvar344[(1'h0):(1'h0)] ?
                      {(wire350 * wire331)} : reg399[(4'h9):(2'h3)]),
                  (^~$unsigned({forvar335}))});
              reg438 = reg395;
              reg439 = ({(~|(reg391 ^~ (reg383 ? reg410 : (8'hb9))))} ?
                  ($signed((wire350 ~^ $signed(forvar421))) >= ($unsigned(wire334) ?
                      reg371 : reg379)) : (|(8'hab)));
              reg440 <= $signed(reg395);
            end
          reg441 = reg351[(1'h1):(1'h0)];
          if ((^reg413[(5'h11):(3'h7)]))
            begin
              reg442 = ((((forvar357 < forvar415) != (&forvar353)) >= (8'ha8)) ?
                  reg382[(1'h1):(1'h1)] : $unsigned($signed({((7'h44) != reg431),
                      reg400})));
              reg443 = ({forvar415,
                  reg397} >> (($unsigned(reg427) ^~ wire327) * (8'ha6)));
              reg444 = reg441;
            end
          else
            begin
              reg442 = {$unsigned((&(~&$unsigned((7'h41)))))};
              reg443 <= (^~$signed($unsigned(forvar390[(4'hd):(2'h3)])));
            end
        end
    end
  assign wire445 = "BbSECRqfUy";
  always
    @(posedge clk) begin
      for (forvar446 = (1'h0); (forvar446 < (1'h0)); forvar446 = (forvar446 + (1'h1)))
        begin
          for (forvar447 = (1'h0); (forvar447 < (2'h2)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 = $unsigned($signed((-reg370)));
              reg449 = ((forvar389[(2'h2):(1'h0)] < $unsigned(reg425[(4'he):(4'ha)])) << $signed(($unsigned((reg412 ?
                  wire445 : forvar426)) << $unsigned({forvar390}))));
              reg450 <= {((reg383[(1'h0):(1'h0)] && reg413) ?
                      reg448 : (^($unsigned(reg373) ^~ ((8'hbd) ?
                          reg379 : (7'h42))))),
                  (|({reg441[(2'h3):(1'h1)], reg386} + {$unsigned(reg382),
                      ((8'ha5) ^~ forvar447)}))};
            end
          for (forvar451 = (1'h0); (forvar451 < (3'h4)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 <= wire401[(3'h7):(3'h6)];
              reg453 <= $unsigned(forvar447);
              reg454 <= ($unsigned("eD8VV") >= (((+reg397) == ($unsigned(wire328) >= (reg352 != reg410))) ?
                  ((~|$signed(reg338)) ?
                      reg367 : reg437) : (~|("" * "2yLIk7CpEnQRO"))));
              reg455 = ((7'h41) ^~ $signed($signed((~&$signed(reg367)))));
            end
          if (reg413)
            begin
              reg456 = (~&forvar372[(4'h8):(1'h1)]);
              reg457 = reg438;
            end
          else
            begin
              reg456 = (-$unsigned(($signed(forvar365) * (8'ha9))));
              reg457 = (((|forvar344) << ($signed((wire332 <= forvar426)) & (~{reg424,
                  reg386}))) <= (^reg370[(1'h0):(1'h0)]));
            end
          reg458 = $unsigned($signed(reg436));
          for (forvar459 = (1'h0); (forvar459 < (1'h1)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 <= $signed($unsigned(((wire445 >= reg450[(2'h3):(1'h0)]) && ((reg428 ?
                  reg373 : (8'hb0)) | reg373[(4'hd):(4'ha)]))));
              reg461 = (forvar357[(2'h3):(1'h0)] ?
                  {$signed((~(reg388 >> reg356))),
                      reg420[(4'ha):(3'h7)]} : reg429);
              reg462 = ($signed((((reg342 >>> wire445) >>> "0LcRai13v8Tz6qhRJdDD") >= (reg352 << reg361))) ?
                  $signed($unsigned(reg423)) : $signed(reg407[(2'h2):(1'h0)]));
              reg463 <= forvar353[(3'h4):(2'h2)];
              reg464 = {reg412[(2'h2):(1'h0)]};
            end
        end
      for (forvar465 = (1'h0); (forvar465 < (3'h4)); forvar465 = (forvar465 + (1'h1)))
        begin
          for (forvar466 = (1'h0); (forvar466 < (1'h1)); forvar466 = (forvar466 + (1'h1)))
            begin
              reg467 = {"wTWUh9Kw4V8q30kArdXg"};
              reg468 = forvar465;
              reg469 <= ($unsigned($unsigned($signed((~|reg413)))) ?
                  reg428[(1'h1):(1'h1)] : (reg347[(1'h1):(1'h0)] ~^ $signed($unsigned($signed(forvar404)))));
              reg470 = forvar430[(3'h5):(3'h4)];
              reg471 <= "FyFT4Ukn";
            end
        end
      reg472 <= ($signed(reg469[(4'h9):(2'h2)]) ?
          (reg406 && ((~|$unsigned((8'hbc))) | $signed($unsigned(reg361)))) : ({($unsigned((8'ha0)) ?
                      $signed(reg410) : $unsigned(reg435)),
                  "k7iHxZalfWX"} ?
              ((reg355[(2'h2):(1'h0)] ?
                  ((8'ha6) ?
                      reg437 : reg409) : $signed(reg458)) ^ $unsigned($signed(reg361))) : reg452));
    end
  assign wire473 = {reg361};
  always
    @(posedge clk) begin
      for (forvar474 = (1'h0); (forvar474 < (1'h1)); forvar474 = (forvar474 + (1'h1)))
        begin
          if (wire330)
            begin
              reg475 <= (((8'h9d) & $signed(forvar364[(2'h2):(2'h2)])) ?
                  (~&$unsigned((^(reg457 ?
                      forvar365 : reg400)))) : $signed(forvar421[(3'h7):(3'h7)]));
              reg476 = (reg347 ?
                  (reg398[(4'he):(4'hd)] || (reg343[(2'h3):(1'h1)] << reg345)) : (forvar364[(1'h1):(1'h1)] ?
                      ($unsigned(reg363[(1'h0):(1'h0)]) >>> (&$unsigned(reg419))) : {reg376[(2'h2):(1'h1)]}));
              reg477 <= (~&(~&($unsigned(reg362[(3'h4):(2'h2)]) ?
                  (reg376 ?
                      reg435[(3'h5):(2'h3)] : forvar446[(2'h2):(2'h2)]) : reg413[(5'h11):(4'hc)])));
              reg478 = (8'ha5);
              reg479 <= (wire473 ^~ reg413[(4'hc):(4'h9)]);
            end
          else
            begin
              reg475 <= (^({reg433,
                  reg362[(2'h3):(2'h3)]} >= $signed((^$unsigned(reg442)))));
              reg476 = $signed((^~($signed($unsigned(reg449)) ?
                  $unsigned((+reg423)) : "Z8")));
            end
          for (forvar480 = (1'h0); (forvar480 < (2'h2)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= $unsigned($signed(reg408));
              reg482 <= {(8'hb1)};
              reg483 <= $unsigned((-(8'h9d)));
            end
          if (($unsigned(reg382) ? reg427 : {reg362}))
            begin
              reg484 = (reg437 ? reg374 : (8'ha0));
              reg485 <= {{reg448[(3'h5):(3'h4)], reg387}};
              reg486 <= "ZMSqDqGZ1cdG0FLlld";
            end
          else
            begin
              reg484 = wire327[(3'h6):(3'h4)];
              reg485 = ($unsigned($signed((8'haf))) ?
                  $unsigned(forvar447[(2'h2):(2'h2)]) : (-reg468[(3'h4):(3'h4)]));
              reg486 <= ($signed(((reg378 | $signed(reg439)) * (!$signed(reg343)))) ?
                  {"FkaplFpNMvuYBoMX"} : (8'ha4));
              reg487 = (7'h42);
            end
        end
      for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
        begin
          reg489 <= {($unsigned((((8'hb1) ? (8'hbb) : reg373) == (forvar446 ?
                  wire401 : reg373))) <= $signed({{wire445, reg416}})),
              (7'h43)};
        end
      for (forvar490 = (1'h0); (forvar490 < (1'h0)); forvar490 = (forvar490 + (1'h1)))
        begin
          reg491 <= $unsigned((|$signed((((8'hb2) ?
              (8'hba) : (8'ha7)) ~^ (^~(8'h9e))))));
          for (forvar492 = (1'h0); (forvar492 < (2'h2)); forvar492 = (forvar492 + (1'h1)))
            begin
              reg493 <= reg481[(4'he):(4'h8)];
              reg494 = $signed(((reg363 | ((~|(8'hbb)) ?
                  (wire445 ?
                      (8'hae) : forvar434) : wire333[(3'h4):(2'h2)])) - forvar421[(3'h7):(3'h4)]));
            end
          for (forvar495 = (1'h0); (forvar495 < (1'h1)); forvar495 = (forvar495 + (1'h1)))
            begin
              reg496 = $unsigned((|("" ?
                  reg399 : $signed(((8'ha6) || forvar417)))));
              reg497 = {(~($unsigned(((8'hae) ^~ reg431)) ?
                      "StW6YSf" : {(forvar446 >> reg379), {(8'ha4)}})),
                  reg470};
              reg498 <= (^~reg494);
              reg499 <= reg423;
            end
          reg500 <= $unsigned((|forvar353));
        end
      for (forvar501 = (1'h0); (forvar501 < (1'h0)); forvar501 = (forvar501 + (1'h1)))
        begin
          reg502 = $unsigned($unsigned($signed(reg487)));
          if ((^~$signed((8'haf))))
            begin
              reg503 = ({(reg362 ? (|(reg479 ? (8'hbd) : reg475)) : (8'hb7)),
                      reg413[(4'h8):(3'h5)]} ?
                  ($signed($signed(((8'ha3) >= reg420))) ?
                      reg469[(1'h1):(1'h0)] : (($signed(reg376) ?
                              $unsigned(reg437) : {forvar344}) ?
                          ((8'h9f) != forvar360) : reg471[(3'h6):(2'h3)])) : (((reg444[(1'h1):(1'h1)] < $signed(wire333)) ?
                      ((reg440 ?
                          (8'hac) : reg497) ~^ (8'hb7)) : $unsigned((reg394 ?
                          reg454 : wire349))) && ((~reg460[(4'ha):(1'h1)]) >> reg398)));
            end
          else
            begin
              reg503 = {$signed({{(~^(8'hb7))}}),
                  (reg393 ?
                      (($unsigned(reg429) ?
                          (-(7'h42)) : $unsigned((8'haa))) <<< reg348[(3'h5):(1'h0)]) : ({(|reg477),
                              $signed(reg433)} ?
                          reg494 : $signed(wire329)))};
              reg504 = $unsigned(reg475);
              reg505 <= {$unsigned({reg370[(1'h1):(1'h1)],
                      $unsigned((reg348 || reg384))})};
              reg506 <= reg343;
              reg507 <= reg484[(1'h0):(1'h0)];
            end
          if ({(8'ha4),
              $unsigned((|((reg387 ? reg370 : (8'hb1)) ?
                  reg475[(2'h3):(2'h2)] : (&reg461))))})
            begin
              reg508 = $unsigned($unsigned($signed(((forvar447 ?
                      forvar501 : (8'ha6)) ?
                  (~^reg497) : (reg369 >>> forvar365)))));
              reg509 <= {reg487[(2'h3):(2'h2)]};
              reg510 <= reg431[(4'h8):(3'h6)];
              reg511 <= reg496;
              reg512 = (~^reg481);
            end
          else
            begin
              reg508 <= reg493[(3'h7):(3'h6)];
            end
          reg513 <= reg469;
          for (forvar514 = (1'h0); (forvar514 < (3'h4)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 <= reg381;
              reg516 = $signed($unsigned($signed(reg438)));
              reg517 = reg384[(4'h9):(3'h4)];
              reg518 <= $signed(((($signed(reg409) ?
                      {reg376} : (reg442 ? reg356 : forvar446)) ?
                  $unsigned($signed(reg424)) : (&(~&(8'hbc)))) && (^~{$signed(reg378),
                  $unsigned((8'hae))})));
              reg519 = ((8'ha9) ?
                  (reg418[(2'h3):(1'h1)] <= $signed(reg369[(2'h2):(1'h0)])) : $unsigned(((reg471 ?
                          $signed(reg462) : reg380) ?
                      {(reg470 ? (8'hb3) : forvar474),
                          (+(8'hb2))} : forvar354[(4'h8):(4'h8)])));
            end
        end
      if (reg512[(2'h3):(2'h3)])
        begin
          for (forvar520 = (1'h0); (forvar520 < (1'h0)); forvar520 = (forvar520 + (1'h1)))
            begin
              reg521 = $unsigned({$signed("CQbt2ni43DCxVCeUH"),
                  reg464[(1'h1):(1'h1)]});
              reg522 <= (~|reg419);
              reg523 <= $unsigned(reg406[(4'ha):(1'h1)]);
            end
        end
      else
        begin
          reg520 <= ((-$signed((~|$signed(reg408)))) ?
              ($signed(reg462) < (reg494 ? reg484 : {{reg380}})) : (((8'hbb) ?
                  $unsigned((-forvar459)) : reg397) | reg370[(3'h4):(1'h0)]));
          for (forvar521 = (1'h0); (forvar521 < (2'h3)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 <= ($signed(forvar346) - $unsigned(reg413[(4'hf):(4'hd)]));
              reg523 <= (~reg428[(1'h0):(1'h0)]);
              reg524 = ((reg414 ?
                      {$signed((wire350 << reg382)),
                          reg457} : ((^~reg374[(4'h9):(2'h3)]) ?
                          $unsigned($signed(reg438)) : (((8'ha0) < reg448) ?
                              $signed(forvar357) : reg498[(3'h4):(2'h3)]))) ?
                  forvar501[(4'h9):(1'h0)] : reg408[(4'he):(3'h6)]);
              reg525 <= (~^{(^reg418[(3'h4):(2'h2)]), {reg523}});
              reg526 = ($unsigned((wire445[(3'h5):(1'h0)] + (reg484 >>> forvar459))) ?
                  (reg517 ?
                      (((forvar446 + reg439) ?
                          $signed(reg513) : (^reg381)) && (reg439[(4'h8):(3'h6)] ?
                          $signed(reg487) : forvar396[(4'hd):(2'h3)])) : (({(8'ha6)} != $unsigned(reg414)) ?
                          $unsigned((reg483 ?
                              reg374 : reg505)) : ($signed(forvar459) ?
                              (reg441 ?
                                  wire350 : reg338) : (reg482 != (8'h9d))))) : "");
            end
          reg527 = reg494;
          for (forvar528 = (1'h0); (forvar528 < (2'h3)); forvar528 = (forvar528 + (1'h1)))
            begin
              reg529 = (reg432[(3'h7):(3'h5)] == reg338[(1'h0):(1'h0)]);
            end
        end
    end
  assign wire530 = reg521;
  assign wire531 = wire327;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module159
#( parameter param323 = {((&(((8'hb0) ~^ (8'hae)) | (+(8'ha8)))) ? (&{((8'hae) >> (8'hb7)), ((8'hb7) ? (7'h42) : (8'hbb))}) : ((7'h40) ? {(^(8'ha5)), ((8'ha2) ? (8'hb5) : (7'h40))} : (((8'h9f) != (7'h42)) ? (~^(7'h40)) : ((8'ha2) ? (8'ha8) : (8'ha9)))))} )
(y, clk, wire163, wire162, wire161, wire160);
  output wire [(32'h6c6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire163;
  input wire [(5'h15):(1'h0)] wire162;
  input wire [(5'h11):(1'h0)] wire161;
  input wire [(5'h11):(1'h0)] wire160;
  wire [(5'h11):(1'h0)] wire322;
  wire signed [(4'h9):(1'h0)] wire321;
  reg signed [(2'h3):(1'h0)] reg320 = (1'h0);
  reg [(5'h14):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg317 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg316 = (1'h0);
  reg [(3'h7):(1'h0)] reg315 = (1'h0);
  reg [(4'ha):(1'h0)] reg314 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg313 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg312 = (1'h0);
  reg [(4'he):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] reg310 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar309 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar308 = (1'h0);
  reg [(4'hb):(1'h0)] reg307 = (1'h0);
  reg signed [(4'he):(1'h0)] reg306 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar305 = (1'h0);
  reg [(5'h14):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar303 = (1'h0);
  reg [(4'ha):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg301 = (1'h0);
  reg [(5'h14):(1'h0)] reg300 = (1'h0);
  reg [(4'h8):(1'h0)] reg299 = (1'h0);
  reg [(3'h4):(1'h0)] reg298 = (1'h0);
  reg [(4'h9):(1'h0)] reg297 = (1'h0);
  reg [(3'h5):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar295 = (1'h0);
  reg [(4'hb):(1'h0)] reg294 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg292 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar291 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg289 = (1'h0);
  reg [(4'hc):(1'h0)] reg288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg287 = (1'h0);
  reg [(5'h10):(1'h0)] reg286 = (1'h0);
  reg [(5'h13):(1'h0)] reg285 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg284 = (1'h0);
  reg [(3'h6):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg282 = (1'h0);
  reg [(4'h9):(1'h0)] forvar281 = (1'h0);
  reg [(4'ha):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg279 = (1'h0);
  reg [(5'h11):(1'h0)] forvar278 = (1'h0);
  reg signed [(4'he):(1'h0)] reg277 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar276 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar273 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar272 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg271 = (1'h0);
  reg [(3'h6):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar263 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar262 = (1'h0);
  wire [(4'hf):(1'h0)] wire261;
  reg [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(3'h4):(1'h0)] reg259 = (1'h0);
  reg [(4'hd):(1'h0)] reg258 = (1'h0);
  reg [(3'h7):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg256 = (1'h0);
  reg signed [(4'he):(1'h0)] reg255 = (1'h0);
  reg [(5'h15):(1'h0)] reg254 = (1'h0);
  reg [(5'h13):(1'h0)] reg253 = (1'h0);
  reg [(4'ha):(1'h0)] reg252 = (1'h0);
  reg [(4'hf):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg250 = (1'h0);
  reg [(2'h3):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg247 = (1'h0);
  reg [(4'h9):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg245 = (1'h0);
  reg [(4'hd):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar243 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg242 = (1'h0);
  reg [(4'hb):(1'h0)] reg241 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg240 = (1'h0);
  reg [(5'h10):(1'h0)] reg239 = (1'h0);
  reg [(4'hb):(1'h0)] reg238 = (1'h0);
  reg [(5'h11):(1'h0)] forvar237 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg236 = (1'h0);
  reg [(3'h5):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg234 = (1'h0);
  reg [(5'h12):(1'h0)] forvar233 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg232 = (1'h0);
  reg [(5'h10):(1'h0)] forvar231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg [(4'hf):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg228 = (1'h0);
  reg [(2'h3):(1'h0)] reg227 = (1'h0);
  reg [(3'h7):(1'h0)] forvar226 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar224 = (1'h0);
  reg [(4'ha):(1'h0)] reg223 = (1'h0);
  reg [(4'hc):(1'h0)] reg222 = (1'h0);
  reg [(2'h2):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg220 = (1'h0);
  reg [(4'hc):(1'h0)] forvar219 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar218 = (1'h0);
  wire signed [(4'he):(1'h0)] wire217;
  wire signed [(4'hb):(1'h0)] wire216;
  reg signed [(4'hc):(1'h0)] reg215 = (1'h0);
  reg [(3'h5):(1'h0)] reg214 = (1'h0);
  reg signed [(4'he):(1'h0)] reg213 = (1'h0);
  reg [(4'ha):(1'h0)] reg212 = (1'h0);
  reg [(2'h3):(1'h0)] reg211 = (1'h0);
  reg [(4'h8):(1'h0)] forvar210 = (1'h0);
  reg [(2'h2):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg208 = (1'h0);
  reg [(5'h10):(1'h0)] reg207 = (1'h0);
  reg [(4'hd):(1'h0)] forvar206 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg205 = (1'h0);
  reg [(4'hf):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg202 = (1'h0);
  reg [(2'h3):(1'h0)] forvar201 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg200 = (1'h0);
  reg [(5'h11):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg197 = (1'h0);
  reg [(4'hf):(1'h0)] reg196 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar195 = (1'h0);
  reg [(4'hb):(1'h0)] forvar194 = (1'h0);
  reg [(4'hb):(1'h0)] reg193 = (1'h0);
  reg [(4'h8):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg191 = (1'h0);
  reg [(2'h3):(1'h0)] reg190 = (1'h0);
  reg [(5'h13):(1'h0)] reg189 = (1'h0);
  reg [(5'h15):(1'h0)] forvar188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(5'h11):(1'h0)] reg186 = (1'h0);
  reg [(4'hb):(1'h0)] reg185 = (1'h0);
  reg [(4'h8):(1'h0)] reg184 = (1'h0);
  reg [(5'h14):(1'h0)] forvar183 = (1'h0);
  reg [(4'he):(1'h0)] forvar182 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg181 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire180;
  wire signed [(2'h3):(1'h0)] wire179;
  wire [(5'h13):(1'h0)] wire178;
  wire [(4'he):(1'h0)] wire177;
  wire signed [(2'h3):(1'h0)] wire176;
  reg signed [(5'h11):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg174 = (1'h0);
  reg [(4'ha):(1'h0)] reg173 = (1'h0);
  reg [(5'h12):(1'h0)] forvar172 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar171 = (1'h0);
  wire [(4'hf):(1'h0)] wire170;
  reg [(3'h4):(1'h0)] reg169 = (1'h0);
  reg [(4'ha):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar167 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar166 = (1'h0);
  reg [(3'h4):(1'h0)] reg165 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire164;
  assign y = {wire322,
                 wire321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 forvar309,
                 forvar308,
                 reg307,
                 reg306,
                 forvar305,
                 reg304,
                 forvar303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 forvar295,
                 reg294,
                 reg293,
                 reg292,
                 forvar291,
                 forvar290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 forvar281,
                 reg280,
                 reg279,
                 forvar278,
                 reg277,
                 forvar276,
                 reg275,
                 reg274,
                 forvar273,
                 forvar272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 forvar262,
                 wire261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 forvar243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 forvar237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 reg232,
                 forvar231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 forvar226,
                 reg225,
                 forvar224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 forvar218,
                 wire217,
                 wire216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 reg209,
                 reg208,
                 reg207,
                 forvar206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 forvar195,
                 forvar194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 forvar188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 forvar183,
                 forvar182,
                 reg181,
                 wire180,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 reg175,
                 reg174,
                 reg173,
                 forvar172,
                 forvar171,
                 wire170,
                 reg169,
                 reg168,
                 forvar167,
                 forvar166,
                 reg165,
                 wire164,
                 (1'h0)};
  assign wire164 = wire162[(5'h11):(3'h5)];
  always
    @(posedge clk) begin
      reg165 = wire161[(3'h7):(3'h6)];
      for (forvar166 = (1'h0); (forvar166 < (2'h3)); forvar166 = (forvar166 + (1'h1)))
        begin
          for (forvar167 = (1'h0); (forvar167 < (1'h1)); forvar167 = (forvar167 + (1'h1)))
            begin
              reg168 = forvar167[(3'h6):(3'h4)];
              reg169 <= (((&$unsigned(reg168)) != (((forvar166 ?
                          wire164 : wire164) ?
                      wire161 : ((8'hb5) || forvar166)) ?
                  (forvar167[(3'h5):(2'h3)] ^ (|wire164)) : $unsigned((wire160 >= reg165)))) == $unsigned(wire162[(4'hb):(3'h5)]));
            end
        end
    end
  assign wire170 = $signed({{(&(~|wire162)), $signed(((8'ha3) >> wire161))},
                       (wire161 ?
                           ("Q" ?
                               $signed(forvar167) : (+forvar167)) : ((^~wire160) ?
                               (wire164 < wire160) : {wire162, reg169}))});
  always
    @(posedge clk) begin
      for (forvar171 = (1'h0); (forvar171 < (1'h1)); forvar171 = (forvar171 + (1'h1)))
        begin
          for (forvar172 = (1'h0); (forvar172 < (2'h3)); forvar172 = (forvar172 + (1'h1)))
            begin
              reg173 = (((((reg165 ? wire164 : reg168) * ((8'hbc) ?
                          wire163 : reg169)) ?
                      wire162 : reg165) - reg165) ?
                  reg165[(1'h1):(1'h1)] : "9JYJ6");
              reg174 <= reg169;
            end
        end
      reg175 = reg169;
    end
  assign wire176 = reg173[(4'h9):(2'h2)];
  assign wire177 = $signed($signed($signed(reg175)));
  assign wire178 = (!$unsigned(reg169[(2'h3):(1'h0)]));
  assign wire179 = (8'haf);
  assign wire180 = $signed(wire177[(3'h4):(1'h1)]);
  always
    @(posedge clk) begin
      reg181 <= wire180;
      for (forvar182 = (1'h0); (forvar182 < (2'h2)); forvar182 = (forvar182 + (1'h1)))
        begin
          for (forvar183 = (1'h0); (forvar183 < (2'h3)); forvar183 = (forvar183 + (1'h1)))
            begin
              reg184 = {(~$signed((((8'hb1) ? reg169 : reg175) ?
                      $signed((8'ha5)) : reg174))),
                  wire160};
              reg185 = wire176[(1'h0):(1'h0)];
              reg186 = $unsigned(wire160[(2'h3):(1'h0)]);
            end
          reg187 = ($unsigned(forvar166[(1'h1):(1'h1)]) ?
              (reg185 ?
                  $signed($signed((forvar166 >= reg168))) : wire176) : (~wire164));
          for (forvar188 = (1'h0); (forvar188 < (2'h2)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= $signed((^~wire176[(1'h0):(1'h0)]));
              reg190 = (({(7'h43)} ?
                      (reg181 <<< ($signed(wire164) ^ (reg186 ^~ wire180))) : (reg168[(4'h8):(2'h2)] <= wire162[(4'ha):(2'h2)])) ?
                  ((($unsigned(wire160) ?
                          {forvar172,
                              reg184} : (~^forvar188)) <<< $unsigned($signed(forvar167))) ?
                      ({$unsigned(reg189),
                          $signed(reg169)} || (wire160[(4'hc):(3'h4)] ?
                          wire178 : wire163[(4'ha):(1'h1)])) : reg174) : (((reg169 ?
                              wire164 : forvar171[(3'h7):(2'h3)]) ?
                          $signed((~^reg181)) : (^~(reg173 | forvar172))) ?
                      $signed(("xE1QI4re" <<< $signed(wire162))) : (^~(~&(8'hb0)))));
              reg191 <= (wire176 ?
                  $unsigned((((wire164 ? wire163 : reg187) ?
                          $unsigned(reg181) : (^~forvar171)) ?
                      forvar172[(4'hf):(3'h6)] : $unsigned((!wire176)))) : {(|reg165[(2'h2):(1'h0)])});
              reg192 <= reg169;
              reg193 <= (~|{$unsigned(((~^(8'h9e)) >> reg185))});
            end
        end
      for (forvar194 = (1'h0); (forvar194 < (2'h3)); forvar194 = (forvar194 + (1'h1)))
        begin
          for (forvar195 = (1'h0); (forvar195 < (2'h2)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 = ((((~$signed(wire160)) ?
                      ((^~reg173) ^~ (wire179 & forvar195)) : $signed(reg173)) - $signed((forvar182 != $unsigned(forvar166)))) ?
                  ({((forvar188 >= reg169) ?
                          reg191 : (reg185 ? wire162 : (8'hb5))),
                      ({(8'ha5), wire179} ?
                          $unsigned(wire176) : $signed(reg168))} >> wire160) : (~|(+reg185)));
              reg197 <= forvar167;
              reg198 = forvar188[(4'hc):(4'ha)];
              reg199 <= reg189[(5'h10):(4'he)];
              reg200 <= $unsigned($signed($signed(reg192)));
            end
          for (forvar201 = (1'h0); (forvar201 < (2'h2)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 = ((!(~|(wire164 ?
                  ((8'hb9) ?
                      wire180 : (8'hbe)) : (8'haf)))) << ((|$signed($signed((8'ha6)))) ?
                  reg187 : $unsigned($unsigned((|(8'hbf))))));
              reg203 <= "";
              reg204 <= $signed(forvar182[(4'he):(1'h0)]);
              reg205 <= $unsigned((forvar195 + (forvar166 >> $unsigned(wire164))));
            end
        end
      for (forvar206 = (1'h0); (forvar206 < (3'h4)); forvar206 = (forvar206 + (1'h1)))
        begin
          if (forvar172[(3'h5):(2'h3)])
            begin
              reg207 = reg189[(5'h13):(1'h0)];
              reg208 = (~($signed(wire178) > wire170));
              reg209 <= (reg189 * (8'hb2));
            end
          else
            begin
              reg207 = $unsigned((~(^~forvar172[(5'h12):(1'h1)])));
              reg208 = $unsigned(forvar183[(3'h6):(2'h3)]);
              reg209 = (((reg189 ?
                      ("m1" ?
                          {wire178} : (reg190 > forvar182)) : wire177[(1'h1):(1'h0)]) ?
                  (reg173[(4'ha):(4'h8)] ~^ (((8'ha5) ?
                      reg186 : forvar166) == $signed(forvar188))) : $unsigned((~^$signed(reg174)))) <<< (($signed((wire163 == forvar172)) * $signed((forvar206 ?
                      reg165 : wire178))) ?
                  reg200[(1'h0):(1'h0)] : (({wire162, reg200} >> ((8'ha8) ?
                          wire177 : forvar182)) ?
                      wire163 : $signed($signed((8'hb1))))));
            end
          for (forvar210 = (1'h0); (forvar210 < (3'h4)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 = forvar194;
              reg212 <= (~reg204[(4'h9):(3'h7)]);
              reg213 = $unsigned((wire170[(1'h1):(1'h1)] | ((!forvar167) ?
                  reg169 : ($unsigned(forvar183) ?
                      (reg189 ? reg187 : (8'hac)) : wire161[(4'he):(4'hc)]))));
            end
        end
      reg214 <= {$signed($signed(reg185))};
    end
  always
    @(posedge clk) begin
      reg215 <= forvar171;
    end
  assign wire216 = {($unsigned($unsigned($signed(reg190))) && ((-$unsigned(reg213)) ?
                           ($signed(reg204) & (|forvar182)) : ((!forvar194) ?
                               reg208 : reg203[(3'h5):(1'h1)]))),
                       wire164};
  assign wire217 = wire164;
  always
    @(posedge clk) begin
      for (forvar218 = (1'h0); (forvar218 < (3'h4)); forvar218 = (forvar218 + (1'h1)))
        begin
          for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 = reg215[(3'h4):(2'h2)];
              reg221 = wire170[(3'h6):(1'h1)];
              reg222 <= "3OOfhHi9XTy";
              reg223 = (forvar182 >> ((((wire163 ~^ forvar183) | {(8'hab),
                          reg189}) ?
                      (wire163[(3'h4):(1'h1)] <<< forvar166) : $signed((forvar218 ?
                          reg200 : reg212))) ?
                  forvar201 : {((forvar166 ?
                          reg181 : reg209) <<< $unsigned(reg207))}));
            end
          for (forvar224 = (1'h0); (forvar224 < (1'h0)); forvar224 = (forvar224 + (1'h1)))
            begin
              reg225 = $unsigned((^~$unsigned($signed(reg184[(1'h0):(1'h0)]))));
            end
          for (forvar226 = (1'h0); (forvar226 < (2'h3)); forvar226 = (forvar226 + (1'h1)))
            begin
              reg227 = {reg199};
              reg228 <= reg223[(3'h7):(1'h1)];
            end
          reg229 <= (|reg227);
          reg230 <= {(+reg221[(2'h2):(1'h1)]), reg229[(4'hd):(3'h4)]};
        end
    end
  always
    @(posedge clk) begin
      for (forvar231 = (1'h0); (forvar231 < (1'h0)); forvar231 = (forvar231 + (1'h1)))
        begin
          reg232 = {reg220[(1'h1):(1'h1)]};
          for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 <= "IZ1NFubiq60I";
              reg235 <= $unsigned(reg181);
            end
          reg236 = $signed(forvar167);
        end
      for (forvar237 = (1'h0); (forvar237 < (2'h3)); forvar237 = (forvar237 + (1'h1)))
        begin
          reg238 <= (~&({($unsigned(reg214) ?
                  $unsigned(forvar183) : (-reg228))} ^ "XRFt"));
          if ({((((forvar166 << reg211) ? (~^reg199) : reg208) ?
                  $unsigned(reg235) : $unsigned((~&(8'ha1)))) && (^~(~&(forvar194 ^ (8'haf))))),
              ((+("8gDRDJSX3" <<< (&reg174))) ?
                  $signed(((reg232 < (8'hbc)) ?
                      (reg184 ?
                          forvar218 : forvar237) : wire162)) : reg208[(2'h3):(2'h3)])})
            begin
              reg239 = $unsigned($signed(reg168[(1'h1):(1'h0)]));
              reg240 = (8'ha6);
            end
          else
            begin
              reg239 <= reg240;
              reg240 = reg238[(4'hb):(3'h7)];
              reg241 = (!(+(~wire180)));
              reg242 = reg234;
            end
          for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
            begin
              reg244 <= {{{reg174},
                      (reg196 ?
                          ({forvar172, forvar166} >= (reg169 ?
                              wire162 : reg196)) : "8cTN8sQMnHXtU3LIn")}};
              reg245 = $unsigned(forvar237);
              reg246 <= forvar171[(1'h1):(1'h0)];
              reg247 = $unsigned((({$signed(reg242), (~^(8'h9d))} + (+(reg211 ?
                  (8'hba) : forvar226))) + $unsigned($signed(reg236))));
              reg248 <= forvar166[(1'h0):(1'h0)];
            end
          if (($signed({"GMtMiJRWd",
              "h"}) <<< $unsigned((^~{$unsigned(wire177)}))))
            begin
              reg249 <= reg248;
              reg250 <= reg204[(4'hd):(2'h2)];
              reg251 = forvar172[(3'h5):(3'h4)];
            end
          else
            begin
              reg249 <= $signed($unsigned(reg187));
              reg250 <= (wire216 ?
                  forvar206 : (($signed(reg181[(1'h0):(1'h0)]) ?
                      (&reg225) : (~|$signed(wire217))) >= $signed("Sn5mObJnXMpQu")));
              reg251 <= reg203[(1'h0):(1'h0)];
              reg252 = reg242[(4'hc):(3'h4)];
              reg253 = {(((7'h43) > (!$unsigned(reg205))) ?
                      $unsigned($signed((^reg212))) : reg225[(3'h6):(3'h6)])};
            end
          reg254 = "5MBQUK9TLi4GFFa";
        end
      if (reg192)
        begin
          if ("EuhMYrEOUoV6V")
            begin
              reg255 <= (((^~reg208[(2'h2):(1'h1)]) ?
                      reg220[(2'h3):(2'h2)] : (reg207 ?
                          (wire177[(4'hd):(4'h8)] >>> (forvar231 ?
                              reg181 : forvar219)) : reg248)) ?
                  forvar226[(2'h3):(1'h1)] : $signed($signed(reg203)));
              reg256 = $unsigned(((+wire177) != forvar166));
              reg257 <= (!(8'ha4));
              reg258 <= {$unsigned(((((8'hbf) << (8'hbe)) << reg181) * $unsigned("")))};
              reg259 <= reg230;
            end
          else
            begin
              reg255 = $signed((^~reg251));
              reg256 <= {{(!$signed(wire162[(1'h0):(1'h0)])),
                      $signed($unsigned({forvar188, reg208}))},
                  (((((8'haa) ?
                          wire216 : reg203) != {reg222}) == (reg198[(3'h4):(2'h2)] > {reg225})) ?
                      $signed(((reg238 ? reg244 : (8'hbb)) ?
                          (wire164 != reg168) : reg244[(4'ha):(2'h2)])) : ((^(-(7'h41))) + ($signed(reg232) ?
                          $unsigned(wire176) : forvar172[(5'h12):(4'h8)])))};
              reg257 <= {reg175[(4'h8):(3'h4)]};
              reg258 <= reg253[(4'h8):(1'h0)];
            end
          reg260 = reg213;
        end
      else
        begin
          reg255 <= ($signed((8'h9f)) && (forvar243 - wire164));
          reg256 = reg239[(3'h4):(3'h4)];
        end
    end
  assign wire261 = $signed(wire162);
  always
    @(posedge clk) begin
      for (forvar262 = (1'h0); (forvar262 < (2'h2)); forvar262 = (forvar262 + (1'h1)))
        begin
          for (forvar263 = (1'h0); (forvar263 < (2'h2)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 = $unsigned(reg190);
              reg265 <= reg184;
            end
          if (reg223)
            begin
              reg266 = (((~|$unsigned((8'hb8))) ?
                  (~(7'h44)) : $unsigned(reg247[(2'h2):(1'h1)])) || $unsigned(($unsigned($signed((8'hb0))) || $unsigned(wire176))));
              reg267 <= ($signed($signed(reg198)) ?
                  $unsigned(reg221) : $signed((((+reg213) ?
                          (~&forvar263) : (~|wire170)) ?
                      (((7'h43) == reg196) >>> (reg200 || (7'h42))) : reg254)));
              reg268 = $unsigned(forvar171[(3'h6):(3'h6)]);
              reg269 <= (&reg209[(1'h0):(1'h0)]);
              reg270 = (("GmtMNQfftSN6Fz" | reg193) ^ wire170[(2'h3):(2'h3)]);
            end
          else
            begin
              reg266 = $signed($unsigned(($signed($signed(reg229)) ?
                  $unsigned($signed(wire164)) : ((reg208 ? reg268 : reg185) ?
                      wire216 : (forvar237 <<< reg249)))));
            end
          reg271 = {$unsigned(wire170[(4'hf):(4'h9)])};
        end
      for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
        begin
          for (forvar273 = (1'h0); (forvar273 < (3'h4)); forvar273 = (forvar273 + (1'h1)))
            begin
              reg274 = reg271[(4'h8):(3'h6)];
              reg275 = $unsigned($unsigned(reg238[(4'hb):(3'h7)]));
            end
        end
      for (forvar276 = (1'h0); (forvar276 < (2'h2)); forvar276 = (forvar276 + (1'h1)))
        begin
          reg277 = reg220[(3'h6):(3'h5)];
          for (forvar278 = (1'h0); (forvar278 < (2'h3)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= $unsigned(((~|reg223[(1'h0):(1'h0)]) | ((^$unsigned(forvar206)) ?
                  ($signed(reg168) < (^reg264)) : reg257)));
              reg280 = (reg248 & $unsigned((reg245[(3'h6):(3'h6)] >> $unsigned($signed(reg228)))));
            end
          for (forvar281 = (1'h0); (forvar281 < (1'h0)); forvar281 = (forvar281 + (1'h1)))
            begin
              reg282 = (~|"AVwmGynrN");
              reg283 <= {($unsigned({(reg192 | reg214),
                      $unsigned(wire217)}) << (($unsigned(forvar172) - "YH0") > $signed($signed((8'h9c))))),
                  (-$signed(reg253))};
              reg284 = {(((~|(8'hb2)) ^ wire261) << forvar224[(4'hb):(4'h9)])};
            end
          if ({reg202,
              {forvar233,
                  ((~&reg284) ?
                      forvar206 : (reg248 ?
                          ((7'h44) + wire170) : (~^forvar237)))}})
            begin
              reg285 = (forvar262 * $unsigned((~reg277[(3'h6):(2'h2)])));
              reg286 <= "5";
              reg287 = ($signed((+((~^reg220) ?
                  (reg211 * forvar206) : $unsigned(forvar276)))) == $signed(((!((8'hae) ?
                  forvar172 : reg204)) & (forvar262[(4'ha):(3'h5)] ?
                  (7'h44) : forvar188[(5'h11):(4'hf)]))));
            end
          else
            begin
              reg285 <= (|($unsigned($unsigned({reg258})) == forvar206[(4'hd):(1'h1)]));
              reg286 = $signed({{reg193[(4'h8):(1'h1)],
                      {"FqH8QcIFDYL6POAPo", reg260}}});
              reg287 = $signed($signed("oYtTaDNBxnu"));
              reg288 <= $signed(("50R6no3" ^ $unsigned((^(wire180 ?
                  reg265 : reg192)))));
            end
        end
      reg289 = $unsigned(wire164);
      for (forvar290 = (1'h0); (forvar290 < (2'h3)); forvar290 = (forvar290 + (1'h1)))
        begin
          for (forvar291 = (1'h0); (forvar291 < (2'h2)); forvar291 = (forvar291 + (1'h1)))
            begin
              reg292 = (~|wire160[(3'h7):(3'h7)]);
              reg293 <= {(+$signed($signed((reg258 ? forvar167 : reg213)))),
                  $unsigned(forvar195[(1'h1):(1'h1)])};
            end
          reg294 = $signed((&reg275[(4'hb):(3'h7)]));
          for (forvar295 = (1'h0); (forvar295 < (2'h2)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 = $unsigned($signed((8'hb2)));
              reg297 = (!reg191[(3'h4):(2'h3)]);
              reg298 = $unsigned(reg235[(3'h5):(2'h2)]);
            end
          if (($signed(($unsigned(reg292) ?
                  {reg283[(1'h1):(1'h0)],
                      reg229[(4'h9):(4'h8)]} : ($signed(wire161) ?
                      $unsigned(wire163) : (reg294 && (8'hab))))) ?
              reg260 : {{"us2fI0otct7TQWPpV", reg256[(5'h14):(1'h1)]}}))
            begin
              reg299 <= wire180;
              reg300 = $signed({$unsigned((reg259[(1'h0):(1'h0)] ?
                      ((8'ha7) > forvar166) : (reg204 ? reg240 : (8'hac)))),
                  $signed(reg208)});
            end
          else
            begin
              reg299 = "ICKdNwwohrPw0L";
              reg300 <= $signed(reg175);
              reg301 = forvar290;
            end
          reg302 = $unsigned(wire161[(2'h3):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar303 = (1'h0); (forvar303 < (2'h2)); forvar303 = (forvar303 + (1'h1)))
        begin
          reg304 = reg212;
          for (forvar305 = (1'h0); (forvar305 < (1'h1)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 <= reg277[(4'hb):(4'ha)];
              reg307 <= (8'ha7);
            end
        end
      for (forvar308 = (1'h0); (forvar308 < (2'h3)); forvar308 = (forvar308 + (1'h1)))
        begin
          for (forvar309 = (1'h0); (forvar309 < (1'h0)); forvar309 = (forvar309 + (1'h1)))
            begin
              reg310 <= ({$unsigned($signed((reg236 ? (8'hb7) : wire216)))} ?
                  ($signed(reg297) ?
                      ((reg165[(3'h4):(1'h0)] ^ ((8'hba) | reg165)) || (forvar194[(4'h9):(1'h0)] >> (+(8'ha2)))) : reg174[(1'h0):(1'h0)]) : (&reg213));
              reg311 = (reg208 + reg298[(3'h4):(1'h1)]);
            end
          if ({$unsigned($signed(($signed(forvar237) ^~ (~&forvar276))))})
            begin
              reg312 = (~^$unsigned(((reg169 ^~ {reg285, forvar278}) ?
                  (reg246 >>> reg307) : $signed((reg213 ? reg175 : (8'ha5))))));
              reg313 <= $signed({"q0h38"});
              reg314 <= reg232;
              reg315 = (reg288 >> ($signed({(reg169 ? forvar262 : reg247),
                      (forvar210 << reg204)}) ?
                  (forvar166[(1'h0):(1'h0)] && ((forvar278 ? reg221 : (8'hbf)) ?
                      reg208 : forvar295)) : $signed((8'hab))));
            end
          else
            begin
              reg312 = ((^($signed(forvar278) ?
                  reg208 : ((reg222 ~^ forvar231) ?
                      (reg296 > reg277) : $unsigned((8'hbb))))) - ($signed((|(8'hbf))) ?
                  ((reg203 > (forvar263 < (8'hbc))) || ($unsigned((8'h9c)) != reg307[(3'h5):(2'h2)])) : $unsigned(($signed(reg256) ?
                      $signed(forvar171) : (~&reg315)))));
              reg313 <= $signed($signed({$unsigned((wire179 ?
                      forvar303 : reg225)),
                  reg252}));
            end
          reg316 = $unsigned($unsigned($unsigned({(&reg228)})));
          if (reg313)
            begin
              reg317 <= {(((-{(8'ha4)}) * reg304[(4'h9):(3'h5)]) ?
                      ({$unsigned(forvar295)} ?
                          reg316 : ($signed(reg304) ?
                              $signed(reg252) : {reg265,
                                  reg240})) : $signed(("J" ?
                          $signed(reg286) : $unsigned(reg169)))),
                  ($unsigned({$signed(reg288)}) >> ($signed($signed(reg235)) ?
                      (reg297[(4'h8):(2'h3)] <<< $signed((8'hb8))) : $signed(((8'h9d) ?
                          (8'had) : (8'hab)))))};
              reg318 <= reg215;
              reg319 = (((^(+{reg187})) ?
                      ($unsigned($signed(reg283)) ?
                          reg282[(1'h1):(1'h1)] : reg165[(1'h1):(1'h1)]) : reg235[(1'h0):(1'h0)]) ?
                  {(~reg175)} : wire179[(2'h3):(1'h0)]);
            end
          else
            begin
              reg317 <= (-{forvar226, (!$unsigned(reg259[(3'h4):(2'h2)]))});
              reg318 = {(+(&(+$signed(reg191))))};
            end
          reg320 = $signed(forvar166);
        end
    end
  assign wire321 = forvar195[(2'h2):(2'h2)];
  assign wire322 = (^~(~$unsigned(((+(8'ha0)) || reg289))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module708
#( parameter param808 = ((^~(^((^~(8'hbe)) * {(8'hbd)}))) - {((^((8'hb3) ^ (7'h42))) ? {((8'ha6) ? (8'hbd) : (8'ha1)), ((8'hb8) <<< (8'hb0))} : ({(8'hac)} ? (~^(8'hb1)) : (|(8'h9f)))), ({((8'haa) < (8'h9e)), ((8'hba) ? (8'ha2) : (8'hbc))} != (((8'h9d) ? (8'ha7) : (8'ha0)) ~^ (^~(8'hbd))))}) )
(y, clk, wire713, wire712, wire711, wire710, wire709);
  output wire [(32'h4c5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire713;
  input wire [(2'h2):(1'h0)] wire712;
  input wire [(5'h10):(1'h0)] wire711;
  input wire [(4'h8):(1'h0)] wire710;
  input wire [(5'h12):(1'h0)] wire709;
  wire signed [(5'h13):(1'h0)] wire807;
  wire signed [(5'h15):(1'h0)] wire806;
  reg [(5'h10):(1'h0)] reg805 = (1'h0);
  reg [(4'h9):(1'h0)] reg804 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg803 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar802 = (1'h0);
  wire [(4'h8):(1'h0)] wire801;
  wire [(4'hf):(1'h0)] wire800;
  reg signed [(5'h15):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg798 = (1'h0);
  reg [(4'ha):(1'h0)] reg797 = (1'h0);
  reg [(5'h12):(1'h0)] reg796 = (1'h0);
  reg [(3'h6):(1'h0)] reg795 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar794 = (1'h0);
  reg [(5'h10):(1'h0)] forvar793 = (1'h0);
  reg signed [(4'he):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg791 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg790 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg789 = (1'h0);
  reg [(4'hc):(1'h0)] forvar788 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg787 = (1'h0);
  reg [(3'h7):(1'h0)] reg786 = (1'h0);
  reg [(4'ha):(1'h0)] reg785 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg784 = (1'h0);
  reg [(5'h13):(1'h0)] reg783 = (1'h0);
  reg [(4'h8):(1'h0)] reg782 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg781 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar780 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg779 = (1'h0);
  reg [(5'h15):(1'h0)] reg778 = (1'h0);
  reg signed [(4'he):(1'h0)] reg777 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg776 = (1'h0);
  reg [(3'h4):(1'h0)] forvar775 = (1'h0);
  reg [(5'h14):(1'h0)] reg774 = (1'h0);
  reg [(3'h4):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg772 = (1'h0);
  reg [(5'h12):(1'h0)] reg771 = (1'h0);
  reg [(4'h9):(1'h0)] reg770 = (1'h0);
  reg [(5'h10):(1'h0)] forvar769 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar768 = (1'h0);
  wire [(4'hc):(1'h0)] wire767;
  wire [(5'h10):(1'h0)] wire766;
  reg signed [(5'h14):(1'h0)] reg765 = (1'h0);
  reg signed [(4'he):(1'h0)] reg759 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar758 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg757 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg764 = (1'h0);
  reg [(4'hb):(1'h0)] reg763 = (1'h0);
  reg [(4'ha):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg761 = (1'h0);
  reg [(5'h14):(1'h0)] reg760 = (1'h0);
  reg [(4'hf):(1'h0)] forvar759 = (1'h0);
  reg [(3'h7):(1'h0)] reg758 = (1'h0);
  reg [(5'h11):(1'h0)] forvar757 = (1'h0);
  reg [(4'ha):(1'h0)] reg756 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg755 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg754 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar752 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg751 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg750 = (1'h0);
  reg [(4'h9):(1'h0)] reg749 = (1'h0);
  reg [(2'h3):(1'h0)] reg748 = (1'h0);
  reg [(5'h12):(1'h0)] reg747 = (1'h0);
  reg [(5'h11):(1'h0)] forvar746 = (1'h0);
  reg [(3'h5):(1'h0)] reg745 = (1'h0);
  reg [(4'hb):(1'h0)] reg744 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg743 = (1'h0);
  reg [(5'h10):(1'h0)] reg742 = (1'h0);
  reg [(5'h14):(1'h0)] reg741 = (1'h0);
  reg [(4'h8):(1'h0)] forvar740 = (1'h0);
  reg [(3'h6):(1'h0)] forvar739 = (1'h0);
  reg [(2'h3):(1'h0)] reg738 = (1'h0);
  reg [(4'hd):(1'h0)] reg737 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg736 = (1'h0);
  reg [(4'ha):(1'h0)] reg735 = (1'h0);
  reg [(4'h8):(1'h0)] reg734 = (1'h0);
  reg [(3'h6):(1'h0)] reg733 = (1'h0);
  reg [(5'h15):(1'h0)] reg732 = (1'h0);
  reg [(2'h2):(1'h0)] reg731 = (1'h0);
  reg [(5'h13):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'he):(1'h0)] reg729 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg728 = (1'h0);
  reg [(5'h15):(1'h0)] reg727 = (1'h0);
  reg [(5'h14):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar725 = (1'h0);
  reg [(5'h14):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar723 = (1'h0);
  wire [(3'h7):(1'h0)] wire722;
  reg [(5'h14):(1'h0)] reg721 = (1'h0);
  reg [(3'h7):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg719 = (1'h0);
  reg [(5'h14):(1'h0)] reg718 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg717 = (1'h0);
  reg [(4'hc):(1'h0)] forvar716 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar715 = (1'h0);
  wire [(4'ha):(1'h0)] wire714;
  assign y = {wire807,
                 wire806,
                 reg805,
                 reg804,
                 reg803,
                 forvar802,
                 wire801,
                 wire800,
                 reg799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 forvar794,
                 forvar793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 forvar788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 forvar780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 forvar775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 forvar769,
                 forvar768,
                 wire767,
                 wire766,
                 reg765,
                 reg759,
                 forvar758,
                 reg757,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg760,
                 forvar759,
                 reg758,
                 forvar757,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 forvar752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 forvar746,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 forvar740,
                 forvar739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 forvar730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 forvar725,
                 reg724,
                 forvar723,
                 wire722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 forvar716,
                 forvar715,
                 wire714,
                 (1'h0)};
  assign wire714 = ($signed(wire711[(3'h7):(3'h5)]) + $unsigned(($signed(wire710) ^ {{wire713},
                       wire712[(2'h2):(1'h0)]})));
  always
    @(posedge clk) begin
      for (forvar715 = (1'h0); (forvar715 < (3'h4)); forvar715 = (forvar715 + (1'h1)))
        begin
          for (forvar716 = (1'h0); (forvar716 < (2'h3)); forvar716 = (forvar716 + (1'h1)))
            begin
              reg717 <= wire711;
              reg718 <= forvar715[(1'h0):(1'h0)];
              reg719 = $unsigned($signed((((+wire714) ?
                  $signed(forvar716) : "X2X1JzF4ueK") >>> (8'hb5))));
              reg720 = wire712[(1'h0):(1'h0)];
              reg721 = wire713[(4'hc):(4'h8)];
            end
        end
    end
  assign wire722 = $signed(($signed(($signed(wire709) < forvar715)) ?
                       (~^((wire709 || reg720) ?
                           $unsigned(wire714) : (wire710 ?
                               reg720 : reg720))) : {{"qR3e0tmgdop7oB6vE"},
                           wire713[(4'hd):(3'h5)]}));
  always
    @(posedge clk) begin
      for (forvar723 = (1'h0); (forvar723 < (1'h1)); forvar723 = (forvar723 + (1'h1)))
        begin
          if (wire713)
            begin
              reg724 <= reg721;
            end
          else
            begin
              reg724 <= reg724;
            end
          for (forvar725 = (1'h0); (forvar725 < (3'h4)); forvar725 = (forvar725 + (1'h1)))
            begin
              reg726 <= (($unsigned(reg720) ?
                      $signed(({reg724,
                          wire712} - (reg718 ^ (8'haa)))) : ((~^wire714) <= (reg720[(3'h6):(3'h6)] < {forvar716}))) ?
                  $signed(((~&wire711[(1'h1):(1'h0)]) ?
                      ((wire709 ? (8'hb8) : reg717) ?
                          {forvar723, forvar723} : (~&forvar723)) : (|(reg720 ?
                          reg718 : (8'ha5))))) : $signed(((-$signed(reg718)) ?
                      (((8'ha6) ? forvar716 : wire713) ?
                          (^~reg717) : (forvar725 <= reg720)) : $unsigned((forvar716 ?
                          forvar716 : reg719)))));
              reg727 <= ("aGaCFr85v6dDLBOEk" | ((8'hb0) ?
                  $signed($unsigned(forvar716[(3'h4):(3'h4)])) : wire713[(3'h6):(3'h6)]));
              reg728 <= $signed({forvar715});
              reg729 <= forvar725;
            end
          for (forvar730 = (1'h0); (forvar730 < (2'h3)); forvar730 = (forvar730 + (1'h1)))
            begin
              reg731 <= $signed((~reg717));
              reg732 <= (((-$unsigned((reg728 >= forvar716))) <<< $signed(((~^wire722) ?
                      {forvar716, reg720} : (-reg729)))) ?
                  $unsigned(forvar715) : $unsigned((~&reg719)));
              reg733 <= reg717;
              reg734 <= (!(-($signed(((8'hb6) >= reg729)) | $signed((forvar725 <= (8'ha7))))));
            end
          if ($unsigned(($unsigned((^{wire712, wire714})) + ($signed("Pi9MM") ?
              (~&$signed(forvar716)) : ($signed(reg720) ?
                  (wire712 && reg727) : (wire709 ? forvar730 : (8'had)))))))
            begin
              reg735 = (($signed(((wire714 >> forvar716) ?
                          (reg721 ? reg734 : reg720) : (~|(8'h9e)))) ?
                      $unsigned((forvar723 ?
                          wire711[(4'he):(4'h8)] : $signed(reg729))) : $unsigned((!forvar715[(2'h3):(2'h3)]))) ?
                  reg733 : $unsigned((+wire722)));
              reg736 <= reg735[(2'h2):(1'h1)];
              reg737 <= $unsigned((^(forvar730[(5'h11):(4'hd)] - $unsigned((reg728 ?
                  reg727 : wire713)))));
              reg738 <= $unsigned(({reg731[(2'h2):(2'h2)]} | (-((reg733 ?
                      (8'hbd) : (8'ha3)) ?
                  (wire709 || forvar715) : $unsigned(reg735)))));
            end
          else
            begin
              reg735 <= {((({forvar723} & $unsigned(reg724)) ?
                          "IsC6cq3q" : $signed(wire714)) ?
                      ((reg732[(3'h5):(1'h0)] ?
                              (reg729 ?
                                  reg737 : forvar725) : reg738[(2'h2):(1'h0)]) ?
                          wire711[(1'h0):(1'h0)] : $signed((~wire711))) : $unsigned($unsigned((reg732 <<< (8'h9e))))),
                  $unsigned($unsigned($signed((forvar723 + reg729))))};
            end
        end
      for (forvar739 = (1'h0); (forvar739 < (3'h4)); forvar739 = (forvar739 + (1'h1)))
        begin
          for (forvar740 = (1'h0); (forvar740 < (2'h3)); forvar740 = (forvar740 + (1'h1)))
            begin
              reg741 <= wire711;
              reg742 <= ((forvar715[(2'h3):(1'h1)] ~^ reg736[(1'h0):(1'h0)]) - ((~|($signed(wire709) | reg736)) ?
                  {((8'hae) ? $unsigned(forvar723) : (+reg732)),
                      (-$unsigned(wire714))} : forvar739[(1'h1):(1'h0)]));
              reg743 <= $unsigned($signed((wire711[(1'h0):(1'h0)] && "SoC61Y3b")));
              reg744 <= $unsigned((~$unsigned(($signed(wire714) == $signed(reg731)))));
              reg745 = ($signed($signed($signed($unsigned(reg732)))) || forvar716[(1'h1):(1'h0)]);
            end
          for (forvar746 = (1'h0); (forvar746 < (3'h4)); forvar746 = (forvar746 + (1'h1)))
            begin
              reg747 = ((-($unsigned(((8'hbf) ?
                  wire713 : reg727)) < (~|(-reg741)))) == ({(((8'hbd) <<< reg733) && (reg737 ?
                          forvar716 : reg720)),
                      ($signed(reg719) ^ forvar723)} ?
                  {reg719, wire712} : ((forvar740[(3'h7):(1'h1)] ?
                          {wire710} : ((8'haa) <<< forvar716)) ?
                      (wire711[(4'hf):(4'hb)] || $unsigned(reg745)) : forvar716[(3'h5):(3'h5)])));
              reg748 <= {wire711[(3'h4):(2'h3)],
                  ({$signed(forvar716[(4'hc):(4'h8)])} ?
                      $unsigned(($unsigned(reg741) != $unsigned(wire714))) : reg728)};
              reg749 <= {$signed(($unsigned($unsigned(reg717)) ?
                      $signed($unsigned(forvar730)) : $signed((reg747 + wire709)))),
                  $unsigned(({reg731} ? ((~|reg747) | (~^reg734)) : reg719))};
              reg750 = (((~^($signed(wire714) ?
                      (&reg726) : $unsigned(reg719))) ~^ reg729) ?
                  $signed(((reg732 ?
                      $unsigned(reg745) : (~|(8'hab))) == (wire722[(1'h0):(1'h0)] >= {reg731}))) : ((-(reg747 ?
                      (reg729 ?
                          reg736 : reg735) : $signed(forvar739))) | $signed($unsigned(reg738[(1'h1):(1'h1)]))));
              reg751 <= (($unsigned($signed($unsigned(forvar746))) <<< reg737) ~^ $signed(($signed(wire714) ?
                  $signed(reg741) : (((8'hab) ?
                      wire713 : forvar716) && (^~reg744)))));
            end
          for (forvar752 = (1'h0); (forvar752 < (2'h3)); forvar752 = (forvar752 + (1'h1)))
            begin
              reg753 <= forvar723[(5'h13):(5'h11)];
              reg754 = $unsigned((~^$unsigned($unsigned(reg717[(1'h1):(1'h1)]))));
              reg755 = ((~^($signed($signed(reg744)) > $signed((8'ha1)))) ~^ (+(|reg731)));
              reg756 <= reg736;
            end
        end
      if ((&(reg756 ?
          (reg737[(4'h8):(2'h3)] ?
              {$signed(wire710),
                  reg729} : ("BOqvVpYRuKyq" && (reg749 ~^ reg741))) : $unsigned("DsYtSr9"))))
        begin
          for (forvar757 = (1'h0); (forvar757 < (2'h2)); forvar757 = (forvar757 + (1'h1)))
            begin
              reg758 <= {$unsigned(reg717[(1'h0):(1'h0)])};
            end
          for (forvar759 = (1'h0); (forvar759 < (1'h0)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 <= $signed(reg741);
              reg761 = ($signed(reg728) <= $unsigned({({(8'hb4), reg733} ?
                      (reg753 ? reg728 : reg729) : {reg744, forvar723})}));
              reg762 <= $unsigned((~^reg732));
              reg763 = $unsigned($signed((($signed(wire711) ?
                      (8'ha2) : (&reg755)) ?
                  (reg732 ?
                      (reg721 >>> (8'hbe)) : (forvar715 ?
                          (8'hae) : reg743)) : forvar725[(3'h4):(3'h4)])));
              reg764 <= $unsigned({$signed(reg749), reg736[(4'ha):(2'h3)]});
            end
        end
      else
        begin
          reg757 = "BdGJCbS";
          for (forvar758 = (1'h0); (forvar758 < (2'h3)); forvar758 = (forvar758 + (1'h1)))
            begin
              reg759 = $signed("xYbuO");
              reg760 <= (({((~|reg764) << (forvar746 ?
                      reg733 : reg751))} <<< $signed((~&forvar752[(4'h9):(3'h4)]))) | $signed(({(reg721 >>> reg728)} >>> (((8'hbb) ?
                      reg757 : reg718) ?
                  {(8'hbd)} : (reg737 ? wire712 : (8'haa))))));
              reg761 = reg744[(4'hb):(4'h9)];
              reg762 <= $unsigned(forvar740[(1'h1):(1'h1)]);
              reg763 <= {"AGqNNGfP"};
            end
        end
      reg765 = ($unsigned($unsigned(reg756[(2'h3):(2'h2)])) ?
          reg734 : "zxL3UlfW4P");
    end
  assign wire766 = wire714;
  assign wire767 = (~^(((forvar740 ?
                           (reg729 || forvar759) : (wire766 ?
                               reg756 : reg750)) ?
                       $signed($unsigned(reg717)) : $unsigned(forvar758)) - ((reg765 ?
                           ((8'hab) != wire709) : "UDz") ?
                       ((forvar730 ?
                           forvar759 : reg762) >= reg750) : $signed($signed(wire710)))));
  always
    @(posedge clk) begin
      for (forvar768 = (1'h0); (forvar768 < (1'h0)); forvar768 = (forvar768 + (1'h1)))
        begin
          for (forvar769 = (1'h0); (forvar769 < (1'h0)); forvar769 = (forvar769 + (1'h1)))
            begin
              reg770 = (~($signed(forvar716[(4'hc):(4'h8)]) ?
                  wire722 : ($unsigned($unsigned((7'h41))) << $unsigned(wire710))));
              reg771 = ((!(forvar739[(3'h5):(2'h2)] ?
                  (((8'hb7) - reg728) ?
                      (reg718 ?
                          (8'hb6) : reg753) : reg726[(2'h3):(2'h2)]) : reg736)) != $signed(reg724[(2'h3):(2'h3)]));
              reg772 = (reg762 ?
                  $signed($signed((+(~&forvar725)))) : ((8'ha8) ?
                      (((~&reg745) - $signed(forvar715)) <<< (^$unsigned(reg743))) : $signed("Z4qgi")));
              reg773 <= (forvar752 ~^ $signed(forvar715[(2'h3):(1'h1)]));
            end
          reg774 <= $unsigned($unsigned((^$signed((-(8'h9d))))));
          for (forvar775 = (1'h0); (forvar775 < (1'h1)); forvar775 = (forvar775 + (1'h1)))
            begin
              reg776 <= (^reg751[(3'h7):(1'h0)]);
              reg777 = $signed(($unsigned(reg771) ?
                  {$unsigned((reg726 ? reg733 : reg759)),
                      $unsigned((reg729 ^ wire766))} : ((~|{wire714,
                      reg745}) ^~ (8'ha8))));
              reg778 <= $signed(reg750);
            end
          reg779 <= "XeI";
        end
      for (forvar780 = (1'h0); (forvar780 < (2'h2)); forvar780 = (forvar780 + (1'h1)))
        begin
          if (reg760)
            begin
              reg781 <= (forvar740[(3'h5):(1'h0)] + {$signed($signed($unsigned(reg717))),
                  $signed($signed((-wire766)))});
              reg782 <= $signed(reg781);
            end
          else
            begin
              reg781 = forvar739[(3'h5):(3'h4)];
              reg782 = reg738;
              reg783 = $unsigned($unsigned(((^~(forvar716 ?
                      forvar757 : reg762)) ?
                  ($unsigned(wire709) & reg743[(4'h8):(3'h7)]) : $unsigned(((8'hbe) ?
                      (8'ha4) : reg757)))));
              reg784 <= $unsigned((reg731[(2'h2):(1'h1)] ?
                  {(7'h44)} : {((forvar780 >= reg773) << (forvar716 ^ reg755))}));
              reg785 <= {($unsigned((!$unsigned(forvar725))) ?
                      ($unsigned($unsigned(reg757)) ?
                          (forvar768[(5'h10):(4'hd)] >> (reg720 ?
                              reg773 : (8'haf))) : $unsigned((forvar758 < reg732))) : reg772[(3'h6):(2'h3)])};
            end
          reg786 = {((!((reg749 >>> reg778) ?
                  $signed(forvar716) : $unsigned((8'hb4)))) != reg738[(2'h2):(1'h0)]),
              (reg782 ?
                  (~&(!$signed(forvar758))) : ((^~(wire711 >>> (8'hb8))) ?
                      reg724[(3'h5):(2'h3)] : wire712[(1'h0):(1'h0)]))};
          reg787 = (($unsigned((-$signed(reg717))) - reg784) ?
              $signed($unsigned((~^(reg718 > reg770)))) : (reg745 != $signed(reg721)));
          for (forvar788 = (1'h0); (forvar788 < (1'h1)); forvar788 = (forvar788 + (1'h1)))
            begin
              reg789 <= $unsigned(forvar715);
              reg790 <= (reg750 & (8'ha9));
              reg791 <= ($signed($unsigned($signed(reg771))) ^~ wire714);
            end
          reg792 = $unsigned($unsigned(forvar769[(4'he):(4'h9)]));
        end
      for (forvar793 = (1'h0); (forvar793 < (1'h1)); forvar793 = (forvar793 + (1'h1)))
        begin
          for (forvar794 = (1'h0); (forvar794 < (2'h2)); forvar794 = (forvar794 + (1'h1)))
            begin
              reg795 = (^~(|(+$signed((forvar793 ? reg727 : reg748)))));
              reg796 <= reg756;
              reg797 = forvar780;
              reg798 <= (|(&(forvar715[(2'h3):(2'h2)] ^ $unsigned((reg795 ?
                  reg787 : reg771)))));
            end
          reg799 = $unsigned(reg754[(2'h3):(1'h0)]);
        end
    end
  assign wire800 = $unsigned($signed((forvar746[(3'h6):(3'h6)] ?
                       reg784 : (-{(8'hb1)}))));
  assign wire801 = (reg731[(1'h0):(1'h0)] ?
                       reg747[(4'ha):(1'h0)] : (&(reg756 || (^~reg785))));
  always
    @(posedge clk) begin
      for (forvar802 = (1'h0); (forvar802 < (1'h1)); forvar802 = (forvar802 + (1'h1)))
        begin
          if ((reg726 & $unsigned((~^{reg777, (~^wire712)}))))
            begin
              reg803 = $unsigned($signed((^$signed((reg757 ?
                  reg737 : forvar780)))));
              reg804 = ($signed(($signed(reg721[(5'h14):(4'h9)]) ?
                      (&forvar775[(1'h0):(1'h0)]) : (8'ha2))) ?
                  (($signed(reg732) | (+(~|forvar802))) > (8'hb8)) : {reg721[(4'hd):(4'hb)],
                      (($unsigned(forvar746) > (wire709 ?
                              forvar757 : forvar730)) ?
                          ((reg795 ? reg771 : reg770) ?
                              $unsigned(reg717) : {forvar725}) : reg726[(5'h13):(4'hd)])});
              reg805 <= ($signed($signed({(reg777 & reg761),
                  (wire800 ?
                      reg757 : forvar758)})) > (~^$signed($unsigned($unsigned((8'h9d))))));
            end
          else
            begin
              reg803 <= reg726;
              reg804 = (reg720 - (8'h9d));
            end
        end
    end
  assign wire806 = ({$unsigned("PuoinxkpOKZSQlr"), reg728[(3'h4):(1'h1)]} ?
                       $unsigned((({(8'h9e), wire712} ^~ ((8'hb8) ?
                           wire712 : forvar802)) != reg734)) : (({$unsigned(reg797)} == (+reg777[(4'hd):(4'h8)])) ?
                           {$unsigned((reg771 ~^ forvar794)),
                               (reg749[(2'h2):(1'h1)] * {(8'hb8)})} : "w6"));
  assign wire807 = (reg753 ^~ (~|$signed((^(reg759 * reg748)))));
endmodule
module top
#(parameter param747 = (8'hb4), parameter param748 = param747)
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h8f1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire0;
  input wire [(5'h12):(1'h0)] wire1;
  input wire signed [(4'hd):(1'h0)] wire2;
  input wire signed [(3'h4):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire4;  
  reg [(5'h13):(1'h0)] reg181 = (1'h0);
  reg signed [(4'he):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg199 = (1'h0);
  reg [(5'h15):(1'h0)] forvar193 = (1'h0);
  assign y = {wire218,
                 wire217,
                 wire216,
                 wire215,
                 (1'h0)};
  assign wire215 = forvar193[(4'hb):(2'h3)];
  assign wire216 = reg199[(2'h3):(2'h3)];
  assign wire217 = (^~reg149);
  assign wire218 = (-reg181[(5'h13):(4'h8)]);
endmodule

module module246  (y, clk, wire247, wire248, wire249, wire250);
  output wire [(32'h3ba):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire247;
  input wire signed [(4'h8):(1'h0)] wire248;
  input wire signed [(5'h11):(1'h0)] wire249;
  input wire signed [(3'h5):(1'h0)] wire250;
  reg [(4'ha):(1'h0)] reg717 = (1'h0);
  reg [(4'he):(1'h0)] reg716 = (1'h0);
  reg [(4'hf):(1'h0)] reg715 = (1'h0);
  reg [(5'h15):(1'h0)] reg714 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg713 = (1'h0);
  reg [(3'h4):(1'h0)] forvar712 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg711 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg709 = (1'h0);
  reg [(2'h3):(1'h0)] reg708 = (1'h0);
  reg [(2'h3):(1'h0)] reg707 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar706 = (1'h0);
  reg [(3'h6):(1'h0)] reg705 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg704 = (1'h0);
  reg [(4'hd):(1'h0)] reg703 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg702 = (1'h0);
  reg [(5'h14):(1'h0)] forvar701 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg700 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg699 = (1'h0);
  reg [(5'h14):(1'h0)] reg698 = (1'h0);
  reg [(4'h9):(1'h0)] forvar697 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg696 = (1'h0);
  reg [(5'h13):(1'h0)] reg695 = (1'h0);
  reg [(5'h10):(1'h0)] forvar694 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg693 = (1'h0);
  reg [(5'h14):(1'h0)] forvar692 = (1'h0);
  reg [(5'h15):(1'h0)] forvar691 = (1'h0);
  wire [(3'h4):(1'h0)] wire689;
  wire [(3'h5):(1'h0)] wire385;
  wire signed [(5'h11):(1'h0)] wire384;
  reg [(4'h9):(1'h0)] forvar251 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg253 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg254 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar256 = (1'h0);
  reg [(3'h6):(1'h0)] reg257 = (1'h0);
  reg [(3'h7):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg260 = (1'h0);
  reg [(4'hc):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar262 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar263 = (1'h0);
  reg [(4'hf):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg265 = (1'h0);
  reg [(4'h8):(1'h0)] reg266 = (1'h0);
  reg signed [(4'he):(1'h0)] reg267 = (1'h0);
  reg [(5'h12):(1'h0)] forvar268 = (1'h0);
  reg [(5'h11):(1'h0)] reg269 = (1'h0);
  reg [(5'h10):(1'h0)] forvar270 = (1'h0);
  reg [(4'hb):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg272 = (1'h0);
  reg [(5'h12):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg275 = (1'h0);
  reg [(5'h11):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar277 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg278 = (1'h0);
  reg [(2'h3):(1'h0)] reg279 = (1'h0);
  reg [(5'h14):(1'h0)] reg280 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg281 = (1'h0);
  reg signed [(4'he):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg283 = (1'h0);
  reg [(4'hb):(1'h0)] reg284 = (1'h0);
  reg [(2'h3):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar286 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar287 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg288 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg290 = (1'h0);
  reg [(4'hb):(1'h0)] reg291 = (1'h0);
  reg [(4'he):(1'h0)] forvar292 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg295 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg297 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire382;
  assign y = {reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 forvar712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 forvar706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 forvar701,
                 reg700,
                 reg699,
                 reg698,
                 forvar697,
                 reg696,
                 reg695,
                 forvar694,
                 reg693,
                 forvar692,
                 forvar691,
                 wire689,
                 wire385,
                 wire384,
                 forvar251,
                 forvar252,
                 reg253,
                 reg254,
                 reg255,
                 forvar256,
                 reg257,
                 reg258,
                 reg259,
                 reg260,
                 reg261,
                 forvar262,
                 forvar263,
                 reg264,
                 reg265,
                 reg266,
                 reg267,
                 forvar268,
                 reg269,
                 forvar270,
                 reg271,
                 reg272,
                 reg273,
                 reg274,
                 reg275,
                 reg276,
                 forvar277,
                 reg278,
                 reg279,
                 reg280,
                 reg281,
                 reg282,
                 reg283,
                 reg284,
                 reg285,
                 forvar286,
                 forvar287,
                 reg288,
                 reg289,
                 reg290,
                 reg291,
                 forvar292,
                 reg293,
                 reg294,
                 reg295,
                 reg296,
                 reg297,
                 wire382,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar251 = (1'h0); (forvar251 < (3'h4)); forvar251 = (forvar251 + (1'h1)))
        begin
          for (forvar252 = (1'h0); (forvar252 < (1'h1)); forvar252 = (forvar252 + (1'h1)))
            begin
              reg253 <= ((~|$unsigned($unsigned((~wire248)))) >> $unsigned(forvar251[(3'h4):(1'h0)]));
              reg254 <= (forvar252[(2'h2):(1'h1)] ?
                  $unsigned($signed((reg253 & $signed(wire248)))) : $unsigned(forvar251[(3'h5):(1'h1)]));
              reg255 = forvar252[(1'h0):(1'h0)];
            end
          for (forvar256 = (1'h0); (forvar256 < (3'h4)); forvar256 = (forvar256 + (1'h1)))
            begin
              reg257 = wire248;
              reg258 <= (reg257[(1'h1):(1'h0)] <= (wire248 ?
                  (~^{((8'had) ? wire248 : (8'hbd)),
                      (wire250 ?
                          wire248 : wire247)}) : wire248[(1'h1):(1'h0)]));
            end
          if ($signed(($unsigned(wire249[(1'h0):(1'h0)]) < reg254[(1'h0):(1'h0)])))
            begin
              reg259 <= (((^{(^wire248), (reg254 < reg255)}) ?
                  $signed($unsigned((wire248 >> wire250))) : (~|$unsigned($unsigned(reg257)))) || $signed("6Ir5szc9fO5"));
              reg260 <= (reg258 ?
                  reg255 : ($signed(($signed(reg258) ?
                          (wire247 <<< reg254) : (^~wire249))) ?
                      $signed(forvar252) : $unsigned({{(7'h44), (8'hbf)},
                          $signed(wire249)})));
              reg261 = $unsigned($signed($signed(reg253[(4'hc):(1'h0)])));
            end
          else
            begin
              reg259 <= (($signed(reg259) >> (~&($signed((8'hab)) ?
                  (forvar251 <= reg253) : $signed(reg257)))) + $signed(($signed({wire249}) && ((|reg260) ?
                  $signed(reg254) : $unsigned((7'h44))))));
              reg260 <= reg255[(2'h3):(1'h1)];
              reg261 <= reg260[(5'h13):(2'h2)];
            end
        end
      for (forvar262 = (1'h0); (forvar262 < (1'h0)); forvar262 = (forvar262 + (1'h1)))
        begin
          for (forvar263 = (1'h0); (forvar263 < (2'h3)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 <= $signed(reg253[(3'h4):(3'h4)]);
              reg265 <= $signed($unsigned({{$signed(reg255)},
                  (((8'hb5) ? forvar252 : reg259) ?
                      (&wire247) : {forvar263, forvar256})}));
              reg266 <= ($unsigned(reg257[(2'h2):(1'h1)]) ?
                  {forvar252[(1'h0):(1'h0)]} : $signed(reg255[(2'h3):(1'h0)]));
            end
          reg267 <= $unsigned($signed($unsigned($unsigned($signed(forvar262)))));
          for (forvar268 = (1'h0); (forvar268 < (1'h1)); forvar268 = (forvar268 + (1'h1)))
            begin
              reg269 <= reg266[(2'h3):(1'h1)];
            end
        end
      for (forvar270 = (1'h0); (forvar270 < (3'h4)); forvar270 = (forvar270 + (1'h1)))
        begin
          if ({(~$unsigned(wire248))})
            begin
              reg271 <= $signed((forvar270[(4'hd):(3'h5)] >= (!reg260[(4'hd):(4'hb)])));
              reg272 <= (~^reg254[(1'h0):(1'h0)]);
              reg273 <= ((reg264[(3'h4):(1'h1)] << {reg266}) ?
                  (forvar252 ?
                      reg253[(4'hc):(2'h2)] : $signed((~&reg260[(5'h11):(2'h3)]))) : $unsigned(((-reg259[(3'h6):(3'h5)]) ?
                      $unsigned(reg255) : wire250)));
              reg274 = reg253[(1'h0):(1'h0)];
            end
          else
            begin
              reg271 = reg267[(4'hb):(1'h0)];
              reg272 <= {(&$signed(((~|forvar270) && "OOaXsZMI3PnY226cISF"))),
                  forvar252};
            end
          if (wire247)
            begin
              reg275 <= (($signed($signed($signed(reg269))) ?
                      (({reg273} ? reg259[(1'h1):(1'h0)] : $signed(wire247)) ?
                          "sKz6didv8iQnJCrkmSNn" : ((reg254 ?
                                  reg272 : wire249) ?
                              (reg267 ~^ reg261) : {reg266})) : wire250[(3'h4):(2'h2)]) ?
                  ("E" ?
                      (~^(~&(7'h44))) : ({reg260[(4'ha):(3'h6)],
                          {wire249}} < $unsigned((forvar251 ?
                          forvar270 : forvar256)))) : $signed((+$signed({reg267,
                      reg261}))));
              reg276 <= reg258;
            end
          else
            begin
              reg275 = $unsigned({$signed(reg259), $signed(reg266)});
            end
          for (forvar277 = (1'h0); (forvar277 < (2'h3)); forvar277 = (forvar277 + (1'h1)))
            begin
              reg278 = reg254;
              reg279 <= $unsigned(forvar251);
              reg280 = ($signed($signed($signed(forvar252))) >> reg260);
              reg281 <= $unsigned($signed($unsigned({reg266})));
              reg282 <= reg260;
            end
          if (reg267)
            begin
              reg283 <= forvar263;
            end
          else
            begin
              reg283 = {$signed($signed(forvar251[(3'h6):(3'h6)]))};
              reg284 <= $signed($unsigned($signed(wire248)));
            end
          reg285 = $signed(reg284[(4'hb):(3'h5)]);
        end
      for (forvar286 = (1'h0); (forvar286 < (3'h4)); forvar286 = (forvar286 + (1'h1)))
        begin
          for (forvar287 = (1'h0); (forvar287 < (2'h3)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 <= $signed((({{wire250, reg260}, wire248} ?
                      "Te0GB3n3" : $signed(((8'haf) ? (8'ha3) : reg264))) ?
                  reg278[(2'h3):(2'h3)] : ("ML5yp" == $signed((reg269 ?
                      forvar263 : reg283)))));
              reg289 = $signed($signed($signed(forvar263)));
              reg290 <= forvar287;
              reg291 <= reg275;
            end
          for (forvar292 = (1'h0); (forvar292 < (3'h4)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 = ((reg260[(1'h0):(1'h0)] != $signed(($signed(reg282) >> forvar268[(1'h1):(1'h0)]))) ?
                  $signed(reg276) : reg273[(4'h9):(1'h0)]);
              reg294 <= {(7'h43), (8'ha4)};
            end
          reg295 <= (&(($signed($signed(forvar277)) - reg273[(4'hd):(3'h7)]) ?
              (reg285 | $signed(reg261[(3'h6):(1'h0)])) : (^~$signed($signed(reg274)))));
          if ($unsigned(reg289))
            begin
              reg296 = reg273[(1'h0):(1'h0)];
              reg297 = (!(-forvar287));
            end
          else
            begin
              reg296 <= $signed(reg297[(1'h1):(1'h0)]);
            end
        end
    end
  assign wire384 = reg261;
  assign wire385 = reg279[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar691 = (1'h0); (forvar691 < (3'h4)); forvar691 = (forvar691 + (1'h1)))
        begin
          for (forvar692 = (1'h0); (forvar692 < (2'h2)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 <= $signed(reg266);
            end
        end
      for (forvar694 = (1'h0); (forvar694 < (3'h4)); forvar694 = (forvar694 + (1'h1)))
        begin
          reg695 = $unsigned(reg282[(4'h9):(3'h7)]);
          reg696 = "VpqP6B2k22WMJuHgWZ";
          for (forvar697 = (1'h0); (forvar697 < (3'h4)); forvar697 = (forvar697 + (1'h1)))
            begin
              reg698 = $unsigned($unsigned(reg260));
              reg699 = $signed({"4iwBauqkC6V6h3",
                  ((8'hbf) ? "9kneuckq0CdONrz" : "K33Kp8mbEE5PIfKSo")});
              reg700 <= reg265;
            end
          for (forvar701 = (1'h0); (forvar701 < (1'h0)); forvar701 = (forvar701 + (1'h1)))
            begin
              reg702 <= $unsigned({reg296[(2'h2):(1'h0)]});
              reg703 <= reg294;
              reg704 <= {$signed(reg290[(3'h6):(2'h2)]),
                  $signed(wire689[(2'h3):(1'h1)])};
              reg705 <= reg258;
            end
        end
      for (forvar706 = (1'h0); (forvar706 < (3'h4)); forvar706 = (forvar706 + (1'h1)))
        begin
          if (reg699[(4'he):(4'he)])
            begin
              reg707 = $signed(((($signed(wire247) ?
                  $unsigned((8'hba)) : (reg257 ?
                      forvar692 : (8'hbb))) || forvar263[(4'ha):(4'ha)]) == (8'h9e)));
              reg708 <= reg260[(4'h8):(3'h7)];
              reg709 <= $unsigned($signed($signed(((|(8'hb9)) ^~ (!reg280)))));
              reg710 = reg259;
              reg711 = {$unsigned(($signed((reg698 ?
                      (8'ha8) : reg710)) != reg700))};
            end
          else
            begin
              reg707 <= ($signed(forvar262[(2'h3):(1'h0)]) >>> $signed({(7'h44),
                  {$unsigned(reg267)}}));
              reg708 <= ($signed((($unsigned(reg257) >= $unsigned((8'ha7))) ?
                      $signed({reg273, reg261}) : ((+forvar286) ?
                          (7'h41) : (-(8'h9c))))) ?
                  forvar270[(2'h3):(1'h0)] : (&$unsigned($signed((+reg291)))));
              reg709 = $unsigned({($unsigned((forvar270 >= reg291)) ?
                      ({reg705} ?
                          (reg279 >> wire247) : forvar287) : {reg258[(2'h2):(1'h1)]}),
                  reg255});
            end
          for (forvar712 = (1'h0); (forvar712 < (1'h0)); forvar712 = (forvar712 + (1'h1)))
            begin
              reg713 = (reg295 ?
                  $signed((^$signed($signed(wire384)))) : reg297);
              reg714 = (~^((^"p3Myzknd3LZD") << wire250[(3'h5):(3'h4)]));
              reg715 <= (reg274[(1'h1):(1'h1)] ?
                  $signed($signed(wire385)) : ($unsigned((|"Lbf0rHmx90HI44")) ?
                      (&reg695) : (((!reg704) ?
                              (reg293 + wire250) : (^forvar287)) ?
                          reg284 : reg294)));
              reg716 <= (|(($signed($unsigned(wire250)) + reg255) ?
                  reg273[(5'h10):(3'h5)] : reg711));
            end
          reg717 = wire382;
        end
    end
endmodule


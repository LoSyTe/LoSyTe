module top
#(parameter param158 = {((8'ha1) + (7'h40))}, parameter param159 = param158)
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h761):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire4;
  input wire signed [(5'h13):(1'h0)] wire3;
  input wire signed [(2'h2):(1'h0)] wire2;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire [(2'h3):(1'h0)] wire0;
  reg [(4'hc):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] reg156 = (1'h0);
  reg [(2'h3):(1'h0)] reg155 = (1'h0);
  reg [(5'h15):(1'h0)] reg154 = (1'h0);
  reg [(4'hf):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg152 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg151 = (1'h0);
  reg [(4'hb):(1'h0)] forvar150 = (1'h0);
  reg [(2'h2):(1'h0)] reg149 = (1'h0);
  reg [(3'h5):(1'h0)] forvar148 = (1'h0);
  reg [(3'h4):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg141 = (1'h0);
  reg [(4'ha):(1'h0)] forvar140 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg146 = (1'h0);
  reg [(4'h9):(1'h0)] reg145 = (1'h0);
  reg [(3'h4):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg142 = (1'h0);
  reg [(2'h2):(1'h0)] forvar141 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg139 = (1'h0);
  reg [(4'he):(1'h0)] reg138 = (1'h0);
  reg [(4'hf):(1'h0)] reg137 = (1'h0);
  reg [(5'h10):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar135 = (1'h0);
  reg [(3'h6):(1'h0)] reg134 = (1'h0);
  reg [(3'h7):(1'h0)] reg133 = (1'h0);
  reg [(4'hb):(1'h0)] reg132 = (1'h0);
  reg [(5'h11):(1'h0)] forvar131 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg130 = (1'h0);
  reg [(5'h12):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg128 = (1'h0);
  reg [(5'h12):(1'h0)] reg127 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar125 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar124 = (1'h0);
  reg [(4'hf):(1'h0)] reg123 = (1'h0);
  reg [(5'h15):(1'h0)] reg122 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg121 = (1'h0);
  reg [(5'h11):(1'h0)] reg120 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg119 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar118 = (1'h0);
  reg [(4'hf):(1'h0)] forvar117 = (1'h0);
  reg [(4'hf):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg115 = (1'h0);
  reg [(5'h14):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg113 = (1'h0);
  reg [(4'hf):(1'h0)] reg112 = (1'h0);
  reg [(5'h11):(1'h0)] forvar111 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar110 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg108 = (1'h0);
  reg [(5'h14):(1'h0)] forvar107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg106 = (1'h0);
  reg [(5'h15):(1'h0)] reg105 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar104 = (1'h0);
  reg [(3'h5):(1'h0)] reg103 = (1'h0);
  reg [(3'h4):(1'h0)] forvar102 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg101 = (1'h0);
  reg [(2'h2):(1'h0)] reg100 = (1'h0);
  reg [(3'h7):(1'h0)] forvar99 = (1'h0);
  reg [(5'h10):(1'h0)] reg98 = (1'h0);
  reg [(4'h8):(1'h0)] forvar97 = (1'h0);
  reg [(5'h10):(1'h0)] forvar96 = (1'h0);
  reg [(5'h12):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg94 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg92 = (1'h0);
  reg [(3'h7):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg90 = (1'h0);
  reg [(5'h12):(1'h0)] reg89 = (1'h0);
  reg [(5'h11):(1'h0)] reg88 = (1'h0);
  reg [(3'h6):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar86 = (1'h0);
  reg [(3'h7):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar84 = (1'h0);
  wire [(4'ha):(1'h0)] wire83;
  reg signed [(2'h3):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(5'h10):(1'h0)] reg80 = (1'h0);
  reg [(4'ha):(1'h0)] reg79 = (1'h0);
  wire [(5'h13):(1'h0)] wire78;
  reg [(4'ha):(1'h0)] reg77 = (1'h0);
  reg [(4'hc):(1'h0)] reg76 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar75 = (1'h0);
  reg [(4'h8):(1'h0)] reg63 = (1'h0);
  reg [(2'h3):(1'h0)] reg74 = (1'h0);
  reg [(2'h2):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg [(3'h5):(1'h0)] forvar70 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg68 = (1'h0);
  reg [(3'h7):(1'h0)] forvar67 = (1'h0);
  reg [(4'h9):(1'h0)] reg66 = (1'h0);
  reg [(5'h15):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg64 = (1'h0);
  reg [(5'h14):(1'h0)] forvar63 = (1'h0);
  reg [(5'h12):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar41 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg40 = (1'h0);
  reg [(4'he):(1'h0)] forvar37 = (1'h0);
  reg [(5'h12):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(4'hf):(1'h0)] reg58 = (1'h0);
  reg [(5'h15):(1'h0)] forvar57 = (1'h0);
  reg [(3'h5):(1'h0)] reg56 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(2'h3):(1'h0)] reg54 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg53 = (1'h0);
  reg [(4'he):(1'h0)] forvar52 = (1'h0);
  reg [(3'h7):(1'h0)] reg51 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar46 = (1'h0);
  reg [(2'h3):(1'h0)] reg45 = (1'h0);
  reg [(3'h5):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg43 = (1'h0);
  reg [(3'h4):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(5'h15):(1'h0)] forvar40 = (1'h0);
  reg [(4'hc):(1'h0)] reg39 = (1'h0);
  reg [(3'h4):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg37 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar35 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg34 = (1'h0);
  reg [(5'h15):(1'h0)] reg33 = (1'h0);
  reg [(3'h7):(1'h0)] reg32 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg30 = (1'h0);
  reg [(5'h10):(1'h0)] forvar29 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg28 = (1'h0);
  reg [(4'hc):(1'h0)] reg27 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg26 = (1'h0);
  reg [(4'ha):(1'h0)] reg25 = (1'h0);
  reg [(3'h5):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar23 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar22 = (1'h0);
  reg [(4'h8):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg20 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg19 = (1'h0);
  reg [(4'h8):(1'h0)] forvar18 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg16 = (1'h0);
  reg [(2'h3):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg [(4'he):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg10 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg12 = (1'h0);
  reg [(4'hd):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar10 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg9 = (1'h0);
  reg signed [(4'he):(1'h0)] reg8 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6 = (1'h0);
  wire [(3'h7):(1'h0)] wire5;
  assign y = {reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 forvar150,
                 reg149,
                 forvar148,
                 reg147,
                 reg141,
                 forvar140,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 forvar141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 reg133,
                 reg132,
                 forvar131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 forvar125,
                 forvar124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 forvar118,
                 forvar117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 forvar111,
                 forvar110,
                 reg109,
                 reg108,
                 forvar107,
                 reg106,
                 reg105,
                 forvar104,
                 reg103,
                 forvar102,
                 reg101,
                 reg100,
                 forvar99,
                 reg98,
                 forvar97,
                 forvar96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 forvar86,
                 reg85,
                 forvar84,
                 wire83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 wire78,
                 reg77,
                 reg76,
                 forvar75,
                 reg63,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 forvar70,
                 reg69,
                 reg68,
                 forvar67,
                 reg66,
                 reg65,
                 reg64,
                 forvar63,
                 reg46,
                 forvar41,
                 reg40,
                 forvar37,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 forvar57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 forvar52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 forvar46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 forvar40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 forvar35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 forvar23,
                 forvar22,
                 reg21,
                 reg20,
                 reg19,
                 forvar18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg10,
                 reg12,
                 reg11,
                 forvar10,
                 reg9,
                 reg8,
                 forvar7,
                 reg6,
                 wire5,
                 (1'h0)};
  assign wire5 = wire1[(5'h11):(2'h2)];
  always
    @(posedge clk) begin
      reg6 <= ((^~($signed({wire2, wire2}) ?
              $unsigned(wire5[(1'h0):(1'h0)]) : wire1)) ?
          wire5[(1'h1):(1'h1)] : wire2[(1'h1):(1'h0)]);
      if (wire5)
        begin
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 <= $signed((-wire1));
            end
          reg9 = $signed($unsigned($unsigned(reg8)));
          for (forvar10 = (1'h0); (forvar10 < (1'h0)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 = $unsigned((-$signed(forvar10[(2'h3):(1'h0)])));
            end
          reg12 <= $unsigned($signed(forvar7));
        end
      else
        begin
          for (forvar7 = (1'h0); (forvar7 < (2'h2)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 <= (7'h40);
              reg9 = wire3;
              reg10 = (wire5[(3'h5):(3'h5)] ?
                  $signed(reg8[(3'h5):(1'h0)]) : reg12);
              reg11 <= ($signed(wire1) ?
                  $signed(wire1) : ((reg10[(5'h12):(4'hd)] ?
                          {((8'ha0) <<< (7'h41))} : "EEHIBr") ?
                      ((~^$unsigned(forvar7)) ?
                          (~|{reg8,
                              (8'ha9)}) : $unsigned((^wire1))) : $unsigned(wire0)));
              reg12 <= ("uHDehs4l8JVaP" >= $signed((8'hb9)));
            end
          reg13 <= reg8[(4'h9):(3'h5)];
          if ($unsigned(($signed($unsigned((wire5 ?
              wire1 : reg6))) ~^ wire1[(4'hd):(2'h3)])))
            begin
              reg14 <= (~|((reg6[(3'h5):(2'h3)] ?
                      (^wire4[(5'h13):(5'h10)]) : ((forvar7 ?
                          (8'hab) : wire1) > wire2)) ?
                  ((^(~reg8)) ?
                      $unsigned($signed(wire1)) : wire5) : ($signed((wire5 ^ (8'hb2))) ?
                      (-$signed(wire0)) : (|((8'ha7) ? wire2 : (8'hb1))))));
            end
          else
            begin
              reg14 = "AbB9r2tS";
              reg15 <= $signed(wire3);
              reg16 = (&($unsigned(reg14) <= {($unsigned(forvar10) ?
                      (wire3 ? wire5 : forvar10) : {(8'ha2)}),
                  ((^reg14) >= $unsigned((8'h9c)))}));
              reg17 <= ({$unsigned((~|reg8)), $unsigned("Q9mF")} > reg11);
            end
          for (forvar18 = (1'h0); (forvar18 < (1'h1)); forvar18 = (forvar18 + (1'h1)))
            begin
              reg19 = ($unsigned(((+wire2[(1'h0):(1'h0)]) ?
                      (&((8'ha1) ? reg17 : reg14)) : {$unsigned(reg8)})) ?
                  $signed(reg11) : (-(~(~^(reg11 >>> forvar7)))));
              reg20 = ($unsigned(($signed((~reg9)) ?
                  reg13[(4'hb):(1'h1)] : wire1[(4'hc):(2'h3)])) <= (&""));
              reg21 <= "CfeHItv7G";
            end
        end
      for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
        begin
          for (forvar23 = (1'h0); (forvar23 < (2'h3)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 <= $signed((|(($unsigned(reg21) ~^ $unsigned(reg13)) ?
                  $signed(reg13) : $signed($unsigned((8'ha3))))));
              reg25 <= forvar7[(2'h2):(1'h0)];
              reg26 = $unsigned($unsigned((reg14[(4'hb):(4'h8)] < $unsigned(reg17))));
              reg27 = (+("7G5XDH" ?
                  (-($signed(reg24) ?
                      reg15[(1'h0):(1'h0)] : (forvar22 ?
                          reg9 : reg10))) : {(-(wire5 >= reg25))}));
              reg28 <= $signed((&$signed(($unsigned((8'hb6)) & (reg9 ?
                  reg13 : wire5)))));
            end
          for (forvar29 = (1'h0); (forvar29 < (3'h4)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 <= $unsigned((~&wire1[(4'hf):(3'h4)]));
              reg31 <= wire1;
            end
          reg32 = wire4;
          reg33 = reg8[(4'hd):(4'ha)];
          reg34 <= (reg13 <<< (($unsigned(((8'hbf) ? reg10 : wire5)) ?
                  (8'hb7) : {(+reg27), (reg6 - reg10)}) ?
              reg15[(1'h0):(1'h0)] : ((+{(8'ha3)}) ?
                  ($signed(reg8) ?
                      reg10 : (reg17 ?
                          reg20 : (7'h42))) : $unsigned(forvar22[(4'hf):(3'h7)]))));
        end
      if ((8'hb2))
        begin
          for (forvar35 = (1'h0); (forvar35 < (2'h2)); forvar35 = (forvar35 + (1'h1)))
            begin
              reg36 <= ({(8'hbd)} ?
                  (reg13[(4'ha):(4'ha)] ^~ $signed($signed($signed((8'ha4))))) : (~&{$unsigned(wire1)}));
              reg37 = reg9[(4'h8):(3'h4)];
              reg38 <= {reg34,
                  ((^((~^wire4) ?
                      ((8'hba) ?
                          reg13 : reg16) : $unsigned(reg30))) != $signed(forvar18))};
              reg39 = $signed($unsigned({$unsigned($signed(reg11)),
                  $signed((+reg37))}));
            end
          for (forvar40 = (1'h0); (forvar40 < (1'h1)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 <= (^~{(reg33[(2'h3):(2'h3)] & "fUdLhnUseUQt3AUCWo")});
              reg42 = $signed($signed($signed(((reg14 || reg30) * forvar7))));
              reg43 <= $unsigned(reg38);
              reg44 <= ($signed("NebLReWdPr2UEQGe") ~^ (|$signed(($unsigned(wire2) <= (reg42 ?
                  (8'hbc) : reg31)))));
              reg45 <= (reg39[(3'h4):(1'h1)] ? $unsigned(reg43) : (7'h41));
            end
          for (forvar46 = (1'h0); (forvar46 < (1'h1)); forvar46 = (forvar46 + (1'h1)))
            begin
              reg47 <= reg15;
              reg48 = (~({{(reg20 ?
                          reg32 : reg10)}} + $unsigned(($signed(reg38) != $unsigned(reg39)))));
              reg49 = reg27[(4'hc):(4'hc)];
              reg50 = ((^reg34) ?
                  $unsigned($signed(($signed(reg27) ^ {reg34,
                      reg12}))) : $signed(($signed($unsigned(reg49)) ?
                      $signed((forvar22 <<< reg42)) : reg41)));
              reg51 <= (~&(($signed(reg43) ?
                  $unsigned($signed(reg9)) : wire2[(1'h0):(1'h0)]) >> $unsigned(($unsigned(reg6) ?
                  $signed(reg44) : {reg30}))));
            end
          for (forvar52 = (1'h0); (forvar52 < (3'h4)); forvar52 = (forvar52 + (1'h1)))
            begin
              reg53 = ($signed(forvar40[(4'h9):(2'h2)]) + reg42[(1'h0):(1'h0)]);
              reg54 <= $unsigned($unsigned($signed($unsigned($unsigned(forvar52)))));
              reg55 <= (8'h9c);
              reg56 = (forvar46[(1'h0):(1'h0)] ? $signed("srlW6iIT") : reg10);
            end
          for (forvar57 = (1'h0); (forvar57 < (2'h2)); forvar57 = (forvar57 + (1'h1)))
            begin
              reg58 <= {(^(!(+$signed(reg28)))),
                  $unsigned((~|(reg8[(2'h2):(1'h1)] ?
                      (^reg10) : reg15[(1'h0):(1'h0)])))};
              reg59 = {{wire1[(4'h9):(4'h9)]}};
              reg60 <= ({($signed(wire2[(1'h0):(1'h0)]) ?
                          (|(~|reg54)) : {((7'h44) ? reg14 : (8'hbb))})} ?
                  $signed(reg10) : forvar18[(1'h1):(1'h0)]);
              reg61 <= $signed(forvar29[(5'h10):(4'hd)]);
              reg62 = reg12;
            end
        end
      else
        begin
          for (forvar35 = (1'h0); (forvar35 < (1'h1)); forvar35 = (forvar35 + (1'h1)))
            begin
              reg36 <= reg54;
            end
          for (forvar37 = (1'h0); (forvar37 < (2'h2)); forvar37 = (forvar37 + (1'h1)))
            begin
              reg38 <= {wire2[(2'h2):(1'h0)]};
              reg39 <= (wire1[(3'h7):(1'h0)] || (8'hbb));
              reg40 <= (~($signed(reg33) <= (($signed(forvar35) ?
                  (forvar46 ?
                      reg16 : reg10) : reg51) || ((8'hac) >>> $unsigned(reg54)))));
            end
          for (forvar41 = (1'h0); (forvar41 < (2'h3)); forvar41 = (forvar41 + (1'h1)))
            begin
              reg42 <= $signed(forvar37[(2'h2):(2'h2)]);
              reg43 <= reg16;
              reg44 <= reg58[(3'h5):(2'h2)];
              reg45 <= "";
              reg46 <= (&(~$unsigned((reg26 * (forvar57 ~^ reg6)))));
            end
          if ($signed(reg26[(1'h1):(1'h1)]))
            begin
              reg47 = ($signed(((8'hbf) ~^ (^(reg53 * forvar7)))) ?
                  {(+($unsigned(reg51) < (+reg60))),
                      reg62[(4'hf):(4'h8)]} : (((|$unsigned(wire2)) << "zmEBNAF5") ?
                      reg34 : $unsigned({(reg10 + (8'haa)), (!reg27)})));
              reg48 <= $unsigned(reg16[(2'h2):(1'h1)]);
              reg49 = ($unsigned(($unsigned(forvar22[(3'h7):(1'h1)]) ?
                      ((forvar57 ? forvar41 : reg53) ?
                          "KNiRH" : (^forvar18)) : $signed($signed(reg20)))) ?
                  reg60[(1'h0):(1'h0)] : $signed((((~^reg59) || forvar10) ?
                      (^(~reg61)) : $signed($signed(reg6)))));
            end
          else
            begin
              reg47 <= $unsigned(((&$signed(reg28)) ?
                  (+(|reg21[(1'h0):(1'h0)])) : forvar10[(2'h3):(1'h1)]));
              reg48 = (^(^{reg50[(3'h4):(2'h3)]}));
            end
          reg50 = (^$unsigned(((((8'haa) ?
              reg30 : reg10) <= reg60) * $unsigned((&reg32)))));
        end
    end
  always
    @(posedge clk) begin
      if (reg34[(4'h9):(1'h1)])
        begin
          for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
            begin
              reg64 <= reg10;
              reg65 <= forvar37;
              reg66 <= $unsigned((($signed(reg40) ^ {reg20}) == (((^(8'hb4)) ?
                      forvar57 : (~&reg50)) ?
                  reg15[(2'h2):(2'h2)] : reg9[(4'hc):(1'h0)])));
            end
          for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= forvar22;
              reg69 <= reg6;
            end
          for (forvar70 = (1'h0); (forvar70 < (1'h1)); forvar70 = (forvar70 + (1'h1)))
            begin
              reg71 <= $unsigned(($unsigned(((^~forvar23) - $signed((8'hb8)))) + ((((8'ha4) && (8'hab)) ?
                  reg48 : forvar57[(3'h4):(2'h3)]) && ((reg66 > reg27) <<< ((8'hbc) ?
                  reg14 : reg20)))));
              reg72 = reg53[(3'h5):(3'h4)];
              reg73 <= (7'h43);
              reg74 <= ({reg46[(3'h7):(3'h5)],
                  ({(reg33 >> forvar70)} <= $signed($unsigned(wire3)))} || reg58);
            end
        end
      else
        begin
          reg63 <= $unsigned(forvar67);
        end
      for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
        begin
          reg76 <= (-("IKdPQMFtEtnoyYmu" + (^~({(8'ha3)} ?
              reg51[(3'h6):(3'h4)] : reg27[(3'h6):(1'h0)]))));
          reg77 <= reg54;
        end
    end
  assign wire78 = "kqYgWCTb9";
  always
    @(posedge clk) begin
      reg79 = (reg47[(3'h5):(3'h4)] ? reg37[(3'h7):(1'h1)] : (7'h43));
      reg80 <= $signed(($signed((!$unsigned(forvar70))) >>> $signed((&(-reg66)))));
      reg81 <= (forvar70[(3'h5):(2'h3)] ?
          (reg59[(2'h3):(2'h3)] >> forvar67[(3'h7):(3'h4)]) : (!$signed(reg55[(3'h4):(2'h2)])));
      reg82 = $signed({$signed(forvar70[(3'h5):(3'h4)])});
    end
  assign wire83 = "5E";
  always
    @(posedge clk) begin
      for (forvar84 = (1'h0); (forvar84 < (3'h4)); forvar84 = (forvar84 + (1'h1)))
        begin
          reg85 <= reg45[(2'h2):(1'h0)];
          for (forvar86 = (1'h0); (forvar86 < (1'h1)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 = reg61;
              reg88 = reg46[(5'h10):(3'h4)];
              reg89 = wire5;
              reg90 <= (-$signed(reg12[(4'h8):(3'h7)]));
              reg91 <= (reg44[(3'h4):(1'h0)] ?
                  ("9H9LyOxUWbMDlRJ5G" ?
                      (($unsigned(forvar37) ?
                              $unsigned((8'h9c)) : reg33[(2'h2):(1'h0)]) ?
                          $signed((!forvar75)) : (wire78[(3'h5):(1'h1)] <= ((8'ha3) ?
                              reg54 : reg64))) : $unsigned(wire5[(3'h6):(2'h2)])) : $signed(($unsigned((+reg21)) <<< forvar46)));
            end
          reg92 <= forvar35;
          if ((&$signed(reg68[(1'h0):(1'h0)])))
            begin
              reg93 <= (({"9DYKiFb",
                  reg74[(2'h3):(1'h1)]} > $signed($unsigned(reg28[(1'h0):(1'h0)]))) ~^ $unsigned($signed((&$unsigned(forvar10)))));
              reg94 = reg72[(2'h3):(1'h1)];
              reg95 <= (forvar52[(4'hb):(2'h2)] != (~&reg32[(3'h7):(3'h5)]));
            end
          else
            begin
              reg93 = (((8'hb2) ^~ (($unsigned((8'hac)) ~^ (reg40 ?
                      reg68 : reg77)) ?
                  reg61 : (reg9 >> ((8'hb3) * reg72)))) >= $signed("4dhODrAb7XTRl"));
              reg94 = (($signed($signed($unsigned(reg48))) ?
                  (~&(!reg56)) : (((reg11 ?
                      forvar52 : (8'hb8)) & (!wire0)) == (&$signed(reg50)))) || (8'ha7));
              reg95 <= reg41;
            end
        end
      for (forvar96 = (1'h0); (forvar96 < (1'h1)); forvar96 = (forvar96 + (1'h1)))
        begin
          for (forvar97 = (1'h0); (forvar97 < (3'h4)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 = (+reg8);
            end
          for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 <= ({reg6, reg68} ?
                  (forvar70 ?
                      (forvar10 ?
                          {(reg62 ?
                                  reg16 : reg61)} : $unsigned((|forvar41))) : reg45) : $unsigned((forvar63[(4'hb):(2'h2)] & $signed(reg61))));
            end
        end
      reg101 = ($unsigned({(reg65 ^ $signed(wire4))}) >> (($signed(((8'ha0) <= (8'haf))) <= forvar10[(1'h1):(1'h0)]) ?
          (&{(forvar75 ?
                  reg24 : forvar46)}) : ($unsigned(reg62[(4'hd):(3'h4)]) ?
              {reg55} : reg6[(4'h9):(3'h4)])));
      for (forvar102 = (1'h0); (forvar102 < (2'h2)); forvar102 = (forvar102 + (1'h1)))
        begin
          reg103 = (((reg45 * $unsigned((~forvar41))) ?
              {$signed((-(8'ha5))),
                  (reg82[(1'h0):(1'h0)] ?
                      reg42 : {reg90,
                          forvar96})} : $unsigned((~$signed(reg90)))) || {(~^(((8'hb2) == forvar96) != $signed(forvar18)))});
          for (forvar104 = (1'h0); (forvar104 < (3'h4)); forvar104 = (forvar104 + (1'h1)))
            begin
              reg105 <= reg92[(3'h4):(1'h1)];
            end
          reg106 <= (reg77 == ((!reg65[(4'hb):(4'hb)]) <<< ($unsigned(reg81) < {"1CPswA7hUzU8hhA",
              $unsigned((8'hac))})));
          for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
            begin
              reg108 = $unsigned(forvar70[(3'h5):(2'h3)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg109 <= $signed((forvar37 ~^ ($signed({reg89, reg49}) ?
          ((forvar57 ? reg90 : reg98) | $signed(reg53)) : $signed((8'hb2)))));
    end
  always
    @(posedge clk) begin
      for (forvar110 = (1'h0); (forvar110 < (1'h1)); forvar110 = (forvar110 + (1'h1)))
        begin
          for (forvar111 = (1'h0); (forvar111 < (2'h3)); forvar111 = (forvar111 + (1'h1)))
            begin
              reg112 <= reg95[(3'h6):(3'h4)];
              reg113 <= (+reg44[(2'h3):(2'h3)]);
              reg114 = (forvar67 ~^ {reg27});
              reg115 <= reg73[(2'h2):(1'h1)];
              reg116 <= $unsigned($signed($unsigned(reg16[(4'hc):(2'h3)])));
            end
        end
      for (forvar117 = (1'h0); (forvar117 < (1'h0)); forvar117 = (forvar117 + (1'h1)))
        begin
          for (forvar118 = (1'h0); (forvar118 < (1'h0)); forvar118 = (forvar118 + (1'h1)))
            begin
              reg119 = $signed((((^~(~|reg6)) << wire4[(3'h4):(2'h3)]) ?
                  (reg61 ?
                      $unsigned((~forvar84)) : ((|reg12) ?
                          reg17[(3'h5):(1'h1)] : $signed(reg32))) : (forvar7 >= ($unsigned(reg71) ?
                      $unsigned(reg115) : (~&forvar23)))));
            end
          if (reg25)
            begin
              reg120 = {($unsigned(((reg24 ? reg19 : (8'hbc)) ?
                          $signed(reg33) : (&reg13))) ?
                      (&reg25[(4'h9):(4'h9)]) : reg115)};
              reg121 <= (reg13[(1'h1):(1'h0)] ^ reg43);
            end
          else
            begin
              reg120 <= (!(((forvar117[(4'h8):(1'h0)] ? {reg31} : reg94) ?
                  (+{(8'ha8),
                      reg120}) : forvar7[(1'h0):(1'h0)]) || {$signed((forvar97 ?
                      forvar67 : forvar37)),
                  wire4[(4'he):(2'h2)]}));
            end
          reg122 <= (~|({forvar40} ~^ $unsigned((forvar75[(3'h7):(3'h4)] ?
              $unsigned(forvar118) : (~&reg71)))));
        end
      reg123 = forvar22[(2'h3):(2'h2)];
      for (forvar124 = (1'h0); (forvar124 < (1'h1)); forvar124 = (forvar124 + (1'h1)))
        begin
          for (forvar125 = (1'h0); (forvar125 < (2'h3)); forvar125 = (forvar125 + (1'h1)))
            begin
              reg126 = $unsigned({$unsigned((^~(reg119 << reg105)))});
              reg127 <= $signed($signed($unsigned(reg79)));
              reg128 = (($signed((((8'hb4) < reg103) ?
                          $unsigned(reg121) : reg28)) ?
                      reg41 : $signed((~(reg11 ? (7'h44) : reg30)))) ?
                  reg8[(4'hc):(4'h9)] : $signed($signed({reg48[(1'h1):(1'h1)]})));
              reg129 = (({$unsigned($unsigned(reg33)),
                  {reg82[(2'h3):(1'h0)],
                      (forvar57 && forvar99)}} <= "mNJTTt") != {(($unsigned((8'ha5)) ?
                          (reg31 && reg76) : ((8'ha5) ^~ reg92)) ?
                      (~&(reg108 ? wire0 : reg109)) : reg115),
                  ("FCw" > $unsigned(reg33[(5'h10):(4'hb)]))});
            end
          reg130 <= (forvar70 ?
              ((((^reg79) ? reg65[(4'hc):(4'h8)] : (~^forvar52)) ?
                  (^~$signed(reg48)) : reg27[(1'h1):(1'h0)]) > $signed($unsigned(forvar10[(3'h5):(3'h4)]))) : {$signed($unsigned((reg85 ?
                      reg12 : forvar96)))});
          for (forvar131 = (1'h0); (forvar131 < (1'h1)); forvar131 = (forvar131 + (1'h1)))
            begin
              reg132 <= ($signed(reg31[(3'h7):(1'h0)]) >>> wire4);
              reg133 <= $unsigned($signed(($unsigned((8'hbd)) < ((~|reg79) <<< reg60[(3'h5):(3'h5)]))));
            end
          reg134 = (!$unsigned((((reg112 ? forvar41 : (8'h9e)) ?
              (reg19 ~^ forvar97) : forvar10[(3'h5):(2'h2)]) > reg81)));
        end
    end
  always
    @(posedge clk) begin
      for (forvar135 = (1'h0); (forvar135 < (1'h0)); forvar135 = (forvar135 + (1'h1)))
        begin
          reg136 = (~|forvar40[(4'hf):(4'ha)]);
          reg137 <= forvar40;
          reg138 = $unsigned(reg16[(3'h4):(3'h4)]);
        end
      reg139 <= (((reg132[(1'h1):(1'h1)] ?
              {(~&reg28), (!reg41)} : ({reg14, (8'hbd)} ?
                  forvar63[(4'ha):(3'h7)] : ((8'ha3) ? reg36 : forvar52))) ?
          (+(((8'hb2) >> reg39) > {(8'hb5), forvar131})) : (8'ha0)) != {{reg27,
              ($signed((7'h40)) ? {forvar84, reg133} : (reg19 > reg59))}});
      if ($unsigned(($unsigned(forvar102[(2'h2):(1'h1)]) ? reg73 : reg134)))
        begin
          reg140 = forvar75;
          for (forvar141 = (1'h0); (forvar141 < (1'h1)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg142 = forvar107;
              reg143 <= reg126;
              reg144 <= wire4[(3'h6):(2'h3)];
              reg145 <= (~reg115);
              reg146 <= (+forvar135);
            end
        end
      else
        begin
          for (forvar140 = (1'h0); (forvar140 < (1'h1)); forvar140 = (forvar140 + (1'h1)))
            begin
              reg141 = (8'h9f);
              reg142 <= {($signed(reg92[(3'h4):(2'h2)]) << reg93), (-forvar67)};
              reg143 = "";
            end
          if ($signed(((($signed(reg14) >>> $unsigned(reg88)) != (forvar131 >>> (~&reg133))) ^ reg146[(4'h9):(3'h4)])))
            begin
              reg144 = reg123[(4'hb):(2'h3)];
            end
          else
            begin
              reg144 <= $signed(($signed((~&(forvar57 ?
                  reg101 : reg119))) ^~ (forvar52[(4'ha):(3'h4)] + $unsigned($unsigned((8'hbf))))));
              reg145 = {(forvar84[(5'h14):(5'h12)] + (((reg142 >= reg38) >>> (+forvar29)) >> ($signed(reg129) * {wire78})))};
              reg146 <= ((^~(-{{wire2, reg85},
                  {forvar140, reg12}})) << reg27[(4'hb):(4'h9)]);
              reg147 = $unsigned(forvar102);
            end
        end
      for (forvar148 = (1'h0); (forvar148 < (1'h1)); forvar148 = (forvar148 + (1'h1)))
        begin
          reg149 <= $unsigned($unsigned(reg142[(1'h0):(1'h0)]));
          for (forvar150 = (1'h0); (forvar150 < (2'h2)); forvar150 = (forvar150 + (1'h1)))
            begin
              reg151 <= {reg61[(3'h7):(1'h1)],
                  (~&($signed(reg49[(1'h0):(1'h0)]) & reg69[(1'h0):(1'h0)]))};
            end
          if (wire2)
            begin
              reg152 <= (reg64[(5'h12):(2'h3)] ?
                  (reg9[(2'h2):(1'h0)] > (8'hba)) : ($unsigned(forvar7[(4'hb):(2'h3)]) ?
                      $signed(reg62[(2'h3):(1'h0)]) : ((-{(8'ha1)}) * forvar7)));
              reg153 = ($unsigned(forvar40[(3'h4):(1'h0)]) > {($unsigned($unsigned(reg15)) && (8'hbe))});
              reg154 = (~&{(-$signed(reg33[(3'h7):(3'h4)]))});
            end
          else
            begin
              reg152 <= (~&$signed(forvar125[(4'ha):(3'h4)]));
              reg153 <= reg6[(4'h8):(3'h4)];
              reg154 = (!{reg74});
              reg155 = $unsigned(($signed(reg90[(3'h7):(3'h4)]) >> ($unsigned(reg100[(1'h1):(1'h1)]) < $unsigned((8'hab)))));
              reg156 = (~|(~^reg119));
            end
        end
      reg157 <= ((~&reg139[(5'h12):(5'h11)]) ?
          $unsigned(($unsigned((reg54 * reg120)) ?
              $signed((~&forvar63)) : "Bg")) : $unsigned(reg48[(5'h14):(4'hc)]));
    end
endmodule